magic
tech sky130A
magscale 1 2
timestamp 1745137735
<< nwell >>
rect -734 178 -312 816
rect 310 -50 732 588
rect 2530 161 2952 214
rect 2530 108 3321 161
rect 2530 37 3690 108
rect 2530 -424 3637 37
rect 2899 -477 3637 -424
rect 3268 -530 3637 -477
rect 4744 -157 5166 -104
rect 4744 -210 5535 -157
rect 4744 -281 5904 -210
rect 4744 -742 5851 -281
rect 5113 -795 5851 -742
rect 5482 -848 5851 -795
rect 6958 -475 7380 -422
rect 6958 -528 7749 -475
rect 6958 -599 8118 -528
rect 6958 -1060 8065 -599
rect 7327 -1113 8065 -1060
rect 7696 -1166 8065 -1113
<< pwell >>
rect -612 -728 -190 92
rect 804 -40 1226 580
rect 1792 249 2214 302
rect 1792 214 2583 249
rect -188 -1086 234 -266
rect 1792 -318 2530 214
rect 2161 -371 2530 -318
rect 3637 -16 4059 37
rect 3637 -69 4428 -16
rect 3637 -104 4797 -69
rect 3637 -583 4744 -104
rect 4006 -636 4744 -583
rect 4375 -689 4744 -636
rect 5851 -334 6273 -281
rect 5851 -387 6642 -334
rect 5851 -422 7011 -387
rect 5851 -901 6958 -422
rect 6220 -954 6958 -901
rect 6589 -1007 6958 -954
rect 8065 -1219 8487 -599
<< nmos >>
rect 1000 170 1030 370
rect -416 -518 -386 -118
rect 1988 -108 2018 92
rect 2357 -161 2387 39
rect 8 -876 38 -476
rect 3833 -373 3863 -173
rect 4202 -426 4232 -226
rect 4571 -479 4601 -279
rect 6047 -691 6077 -491
rect 6416 -744 6446 -544
rect 6785 -797 6815 -597
rect 8261 -1009 8291 -809
<< pmos >>
rect -538 397 -508 597
rect 506 169 536 369
rect 2726 -205 2756 -5
rect 3095 -258 3125 -58
rect 3464 -311 3494 -111
rect 4940 -523 4970 -323
rect 5309 -576 5339 -376
rect 5678 -629 5708 -429
rect 7154 -841 7184 -641
rect 7523 -894 7553 -694
rect 7892 -947 7922 -747
<< ndiff >>
rect 942 358 1000 370
rect 942 182 954 358
rect 988 182 1000 358
rect 942 170 1000 182
rect 1030 358 1088 370
rect 1030 182 1042 358
rect 1076 182 1088 358
rect 1030 170 1088 182
rect -474 -130 -416 -118
rect -474 -506 -462 -130
rect -428 -506 -416 -130
rect -474 -518 -416 -506
rect -386 -130 -328 -118
rect -386 -506 -374 -130
rect -340 -506 -328 -130
rect -386 -518 -328 -506
rect 1930 80 1988 92
rect 1930 -96 1942 80
rect 1976 -96 1988 80
rect 1930 -108 1988 -96
rect 2018 80 2076 92
rect 2018 -96 2030 80
rect 2064 -96 2076 80
rect 2018 -108 2076 -96
rect 2299 27 2357 39
rect 2299 -149 2311 27
rect 2345 -149 2357 27
rect 2299 -161 2357 -149
rect 2387 27 2445 39
rect 2387 -149 2399 27
rect 2433 -149 2445 27
rect 2387 -161 2445 -149
rect -50 -488 8 -476
rect -50 -864 -38 -488
rect -4 -864 8 -488
rect -50 -876 8 -864
rect 38 -488 96 -476
rect 38 -864 50 -488
rect 84 -864 96 -488
rect 38 -876 96 -864
rect 3775 -185 3833 -173
rect 3775 -361 3787 -185
rect 3821 -361 3833 -185
rect 3775 -373 3833 -361
rect 3863 -185 3921 -173
rect 3863 -361 3875 -185
rect 3909 -361 3921 -185
rect 3863 -373 3921 -361
rect 4144 -238 4202 -226
rect 4144 -414 4156 -238
rect 4190 -414 4202 -238
rect 4144 -426 4202 -414
rect 4232 -238 4290 -226
rect 4232 -414 4244 -238
rect 4278 -414 4290 -238
rect 4232 -426 4290 -414
rect 4513 -291 4571 -279
rect 4513 -467 4525 -291
rect 4559 -467 4571 -291
rect 4513 -479 4571 -467
rect 4601 -291 4659 -279
rect 4601 -467 4613 -291
rect 4647 -467 4659 -291
rect 4601 -479 4659 -467
rect 5989 -503 6047 -491
rect 5989 -679 6001 -503
rect 6035 -679 6047 -503
rect 5989 -691 6047 -679
rect 6077 -503 6135 -491
rect 6077 -679 6089 -503
rect 6123 -679 6135 -503
rect 6077 -691 6135 -679
rect 6358 -556 6416 -544
rect 6358 -732 6370 -556
rect 6404 -732 6416 -556
rect 6358 -744 6416 -732
rect 6446 -556 6504 -544
rect 6446 -732 6458 -556
rect 6492 -732 6504 -556
rect 6446 -744 6504 -732
rect 6727 -609 6785 -597
rect 6727 -785 6739 -609
rect 6773 -785 6785 -609
rect 6727 -797 6785 -785
rect 6815 -609 6873 -597
rect 6815 -785 6827 -609
rect 6861 -785 6873 -609
rect 6815 -797 6873 -785
rect 8203 -821 8261 -809
rect 8203 -997 8215 -821
rect 8249 -997 8261 -821
rect 8203 -1009 8261 -997
rect 8291 -821 8349 -809
rect 8291 -997 8303 -821
rect 8337 -997 8349 -821
rect 8291 -1009 8349 -997
<< pdiff >>
rect -596 585 -538 597
rect -596 409 -584 585
rect -550 409 -538 585
rect -596 397 -538 409
rect -508 585 -450 597
rect -508 409 -496 585
rect -462 409 -450 585
rect -508 397 -450 409
rect 448 357 506 369
rect 448 181 460 357
rect 494 181 506 357
rect 448 169 506 181
rect 536 357 594 369
rect 536 181 548 357
rect 582 181 594 357
rect 536 169 594 181
rect 2668 -17 2726 -5
rect 2668 -193 2680 -17
rect 2714 -193 2726 -17
rect 2668 -205 2726 -193
rect 2756 -17 2814 -5
rect 2756 -193 2768 -17
rect 2802 -193 2814 -17
rect 2756 -205 2814 -193
rect 3037 -70 3095 -58
rect 3037 -246 3049 -70
rect 3083 -246 3095 -70
rect 3037 -258 3095 -246
rect 3125 -70 3183 -58
rect 3125 -246 3137 -70
rect 3171 -246 3183 -70
rect 3125 -258 3183 -246
rect 3406 -123 3464 -111
rect 3406 -299 3418 -123
rect 3452 -299 3464 -123
rect 3406 -311 3464 -299
rect 3494 -123 3552 -111
rect 3494 -299 3506 -123
rect 3540 -299 3552 -123
rect 3494 -311 3552 -299
rect 4882 -335 4940 -323
rect 4882 -511 4894 -335
rect 4928 -511 4940 -335
rect 4882 -523 4940 -511
rect 4970 -335 5028 -323
rect 4970 -511 4982 -335
rect 5016 -511 5028 -335
rect 4970 -523 5028 -511
rect 5251 -388 5309 -376
rect 5251 -564 5263 -388
rect 5297 -564 5309 -388
rect 5251 -576 5309 -564
rect 5339 -388 5397 -376
rect 5339 -564 5351 -388
rect 5385 -564 5397 -388
rect 5339 -576 5397 -564
rect 5620 -441 5678 -429
rect 5620 -617 5632 -441
rect 5666 -617 5678 -441
rect 5620 -629 5678 -617
rect 5708 -441 5766 -429
rect 5708 -617 5720 -441
rect 5754 -617 5766 -441
rect 5708 -629 5766 -617
rect 7096 -653 7154 -641
rect 7096 -829 7108 -653
rect 7142 -829 7154 -653
rect 7096 -841 7154 -829
rect 7184 -653 7242 -641
rect 7184 -829 7196 -653
rect 7230 -829 7242 -653
rect 7184 -841 7242 -829
rect 7465 -706 7523 -694
rect 7465 -882 7477 -706
rect 7511 -882 7523 -706
rect 7465 -894 7523 -882
rect 7553 -706 7611 -694
rect 7553 -882 7565 -706
rect 7599 -882 7611 -706
rect 7553 -894 7611 -882
rect 7834 -759 7892 -747
rect 7834 -935 7846 -759
rect 7880 -935 7892 -759
rect 7834 -947 7892 -935
rect 7922 -759 7980 -747
rect 7922 -935 7934 -759
rect 7968 -935 7980 -759
rect 7922 -947 7980 -935
<< ndiffc >>
rect 954 182 988 358
rect 1042 182 1076 358
rect -462 -506 -428 -130
rect -374 -506 -340 -130
rect 1942 -96 1976 80
rect 2030 -96 2064 80
rect 2311 -149 2345 27
rect 2399 -149 2433 27
rect -38 -864 -4 -488
rect 50 -864 84 -488
rect 3787 -361 3821 -185
rect 3875 -361 3909 -185
rect 4156 -414 4190 -238
rect 4244 -414 4278 -238
rect 4525 -467 4559 -291
rect 4613 -467 4647 -291
rect 6001 -679 6035 -503
rect 6089 -679 6123 -503
rect 6370 -732 6404 -556
rect 6458 -732 6492 -556
rect 6739 -785 6773 -609
rect 6827 -785 6861 -609
rect 8215 -997 8249 -821
rect 8303 -997 8337 -821
<< pdiffc >>
rect -584 409 -550 585
rect -496 409 -462 585
rect 460 181 494 357
rect 548 181 582 357
rect 2680 -193 2714 -17
rect 2768 -193 2802 -17
rect 3049 -246 3083 -70
rect 3137 -246 3171 -70
rect 3418 -299 3452 -123
rect 3506 -299 3540 -123
rect 4894 -511 4928 -335
rect 4982 -511 5016 -335
rect 5263 -564 5297 -388
rect 5351 -564 5385 -388
rect 5632 -617 5666 -441
rect 5720 -617 5754 -441
rect 7108 -829 7142 -653
rect 7196 -829 7230 -653
rect 7477 -882 7511 -706
rect 7565 -882 7599 -706
rect 7846 -935 7880 -759
rect 7934 -935 7968 -759
<< psubdiff >>
rect -576 22 -480 56
rect -322 22 -226 56
rect -576 -40 -542 22
rect -260 -40 -226 22
rect 840 510 936 544
rect 1094 510 1190 544
rect 840 448 874 510
rect 1156 448 1190 510
rect 840 30 874 92
rect 1156 30 1190 92
rect 840 -4 936 30
rect 1094 -4 1190 30
rect 1828 232 1924 266
rect 2082 232 2178 266
rect 1828 170 1862 232
rect -576 -658 -542 -596
rect 2144 170 2178 232
rect 1828 -248 1862 -186
rect 2144 -248 2178 -186
rect 1828 -282 1924 -248
rect 2082 -282 2178 -248
rect 2197 179 2293 213
rect 2451 179 2547 213
rect 2197 117 2231 179
rect 2513 117 2547 179
rect 2197 -301 2231 -239
rect 2513 -301 2547 -239
rect -260 -658 -226 -596
rect -576 -692 -480 -658
rect -322 -692 -226 -658
rect -152 -336 -56 -302
rect 102 -336 198 -302
rect 2197 -335 2293 -301
rect 2451 -335 2547 -301
rect -152 -398 -118 -336
rect 164 -398 198 -336
rect -152 -1016 -118 -954
rect 3673 -33 3769 1
rect 3927 -33 4023 1
rect 3673 -95 3707 -33
rect 3989 -95 4023 -33
rect 3673 -513 3707 -451
rect 3989 -513 4023 -451
rect 3673 -547 3769 -513
rect 3927 -547 4023 -513
rect 4042 -86 4138 -52
rect 4296 -86 4392 -52
rect 4042 -148 4076 -86
rect 4358 -148 4392 -86
rect 4042 -566 4076 -504
rect 4358 -566 4392 -504
rect 4042 -600 4138 -566
rect 4296 -600 4392 -566
rect 4411 -139 4507 -105
rect 4665 -139 4761 -105
rect 4411 -201 4445 -139
rect 4727 -201 4761 -139
rect 4411 -619 4445 -557
rect 4727 -619 4761 -557
rect 4411 -653 4507 -619
rect 4665 -653 4761 -619
rect 5887 -351 5983 -317
rect 6141 -351 6237 -317
rect 5887 -413 5921 -351
rect 6203 -413 6237 -351
rect 5887 -831 5921 -769
rect 6203 -831 6237 -769
rect 5887 -865 5983 -831
rect 6141 -865 6237 -831
rect 6256 -404 6352 -370
rect 6510 -404 6606 -370
rect 6256 -466 6290 -404
rect 6572 -466 6606 -404
rect 6256 -884 6290 -822
rect 6572 -884 6606 -822
rect 6256 -918 6352 -884
rect 6510 -918 6606 -884
rect 6625 -457 6721 -423
rect 6879 -457 6975 -423
rect 6625 -519 6659 -457
rect 6941 -519 6975 -457
rect 164 -1016 198 -954
rect 6625 -937 6659 -875
rect 6941 -937 6975 -875
rect 6625 -971 6721 -937
rect 6879 -971 6975 -937
rect -152 -1050 -56 -1016
rect 102 -1050 198 -1016
rect 8101 -669 8197 -635
rect 8355 -669 8451 -635
rect 8101 -731 8135 -669
rect 8417 -731 8451 -669
rect 8101 -1149 8135 -1087
rect 8417 -1149 8451 -1087
rect 8101 -1183 8197 -1149
rect 8355 -1183 8451 -1149
<< nsubdiff >>
rect -698 746 -602 780
rect -444 746 -348 780
rect -698 684 -664 746
rect -382 684 -348 746
rect -698 248 -664 310
rect -382 248 -348 310
rect -698 214 -602 248
rect -444 214 -348 248
rect 346 518 442 552
rect 600 518 696 552
rect 346 456 380 518
rect 662 456 696 518
rect 346 20 380 82
rect 662 20 696 82
rect 346 -14 442 20
rect 600 -14 696 20
rect 2566 144 2662 178
rect 2820 144 2916 178
rect 2566 82 2600 144
rect 2882 82 2916 144
rect 2566 -354 2600 -292
rect 2882 -354 2916 -292
rect 2566 -388 2662 -354
rect 2820 -388 2916 -354
rect 2935 91 3031 125
rect 3189 91 3285 125
rect 2935 29 2969 91
rect 3251 29 3285 91
rect 2935 -407 2969 -345
rect 3251 -407 3285 -345
rect 2935 -441 3031 -407
rect 3189 -441 3285 -407
rect 3304 38 3400 72
rect 3558 38 3654 72
rect 3304 -24 3338 38
rect 3620 -24 3654 38
rect 3304 -460 3338 -398
rect 3620 -460 3654 -398
rect 3304 -494 3400 -460
rect 3558 -494 3654 -460
rect 4780 -174 4876 -140
rect 5034 -174 5130 -140
rect 4780 -236 4814 -174
rect 5096 -236 5130 -174
rect 4780 -672 4814 -610
rect 5096 -672 5130 -610
rect 4780 -706 4876 -672
rect 5034 -706 5130 -672
rect 5149 -227 5245 -193
rect 5403 -227 5499 -193
rect 5149 -289 5183 -227
rect 5465 -289 5499 -227
rect 5149 -725 5183 -663
rect 5465 -725 5499 -663
rect 5149 -759 5245 -725
rect 5403 -759 5499 -725
rect 5518 -280 5614 -246
rect 5772 -280 5868 -246
rect 5518 -342 5552 -280
rect 5834 -342 5868 -280
rect 5518 -778 5552 -716
rect 5834 -778 5868 -716
rect 5518 -812 5614 -778
rect 5772 -812 5868 -778
rect 6994 -492 7090 -458
rect 7248 -492 7344 -458
rect 6994 -554 7028 -492
rect 7310 -554 7344 -492
rect 6994 -990 7028 -928
rect 7310 -990 7344 -928
rect 6994 -1024 7090 -990
rect 7248 -1024 7344 -990
rect 7363 -545 7459 -511
rect 7617 -545 7713 -511
rect 7363 -607 7397 -545
rect 7679 -607 7713 -545
rect 7363 -1043 7397 -981
rect 7679 -1043 7713 -981
rect 7363 -1077 7459 -1043
rect 7617 -1077 7713 -1043
rect 7732 -598 7828 -564
rect 7986 -598 8082 -564
rect 7732 -660 7766 -598
rect 8048 -660 8082 -598
rect 7732 -1096 7766 -1034
rect 8048 -1096 8082 -1034
rect 7732 -1130 7828 -1096
rect 7986 -1130 8082 -1096
<< psubdiffcont >>
rect -480 22 -322 56
rect -576 -596 -542 -40
rect 936 510 1094 544
rect 840 92 874 448
rect 1156 92 1190 448
rect 936 -4 1094 30
rect 1924 232 2082 266
rect -260 -596 -226 -40
rect 1828 -186 1862 170
rect 2144 -186 2178 170
rect 1924 -282 2082 -248
rect 2293 179 2451 213
rect 2197 -239 2231 117
rect 2513 -239 2547 117
rect -480 -692 -322 -658
rect -56 -336 102 -302
rect 2293 -335 2451 -301
rect -152 -954 -118 -398
rect 164 -954 198 -398
rect 3769 -33 3927 1
rect 3673 -451 3707 -95
rect 3989 -451 4023 -95
rect 3769 -547 3927 -513
rect 4138 -86 4296 -52
rect 4042 -504 4076 -148
rect 4358 -504 4392 -148
rect 4138 -600 4296 -566
rect 4507 -139 4665 -105
rect 4411 -557 4445 -201
rect 4727 -557 4761 -201
rect 4507 -653 4665 -619
rect 5983 -351 6141 -317
rect 5887 -769 5921 -413
rect 6203 -769 6237 -413
rect 5983 -865 6141 -831
rect 6352 -404 6510 -370
rect 6256 -822 6290 -466
rect 6572 -822 6606 -466
rect 6352 -918 6510 -884
rect 6721 -457 6879 -423
rect 6625 -875 6659 -519
rect 6941 -875 6975 -519
rect 6721 -971 6879 -937
rect -56 -1050 102 -1016
rect 8197 -669 8355 -635
rect 8101 -1087 8135 -731
rect 8417 -1087 8451 -731
rect 8197 -1183 8355 -1149
<< nsubdiffcont >>
rect -602 746 -444 780
rect -698 310 -664 684
rect -382 310 -348 684
rect -602 214 -444 248
rect 442 518 600 552
rect 346 82 380 456
rect 662 82 696 456
rect 442 -14 600 20
rect 2662 144 2820 178
rect 2566 -292 2600 82
rect 2882 -292 2916 82
rect 2662 -388 2820 -354
rect 3031 91 3189 125
rect 2935 -345 2969 29
rect 3251 -345 3285 29
rect 3031 -441 3189 -407
rect 3400 38 3558 72
rect 3304 -398 3338 -24
rect 3620 -398 3654 -24
rect 3400 -494 3558 -460
rect 4876 -174 5034 -140
rect 4780 -610 4814 -236
rect 5096 -610 5130 -236
rect 4876 -706 5034 -672
rect 5245 -227 5403 -193
rect 5149 -663 5183 -289
rect 5465 -663 5499 -289
rect 5245 -759 5403 -725
rect 5614 -280 5772 -246
rect 5518 -716 5552 -342
rect 5834 -716 5868 -342
rect 5614 -812 5772 -778
rect 7090 -492 7248 -458
rect 6994 -928 7028 -554
rect 7310 -928 7344 -554
rect 7090 -1024 7248 -990
rect 7459 -545 7617 -511
rect 7363 -981 7397 -607
rect 7679 -981 7713 -607
rect 7459 -1077 7617 -1043
rect 7828 -598 7986 -564
rect 7732 -1034 7766 -660
rect 8048 -1034 8082 -660
rect 7828 -1130 7986 -1096
<< poly >>
rect -556 678 -490 694
rect -556 644 -540 678
rect -506 644 -490 678
rect -556 628 -490 644
rect -538 597 -508 628
rect -538 370 -508 397
rect 488 450 554 466
rect 488 416 504 450
rect 538 416 554 450
rect 488 400 554 416
rect 506 369 536 400
rect 506 142 536 169
rect -434 -46 -368 -30
rect -434 -80 -418 -46
rect -384 -80 -368 -46
rect -434 -96 -368 -80
rect 982 442 1048 458
rect 982 408 998 442
rect 1032 408 1048 442
rect 982 392 1048 408
rect 1000 370 1030 392
rect 1000 148 1030 170
rect 982 132 1048 148
rect 982 98 998 132
rect 1032 98 1048 132
rect 982 82 1048 98
rect -416 -118 -386 -96
rect -416 -544 -386 -518
rect 1970 164 2036 180
rect 1970 130 1986 164
rect 2020 130 2036 164
rect 1970 114 2036 130
rect 1988 92 2018 114
rect 1988 -130 2018 -108
rect 1970 -146 2036 -130
rect 1970 -180 1986 -146
rect 2020 -180 2036 -146
rect 1970 -196 2036 -180
rect 2339 111 2405 127
rect 2339 77 2355 111
rect 2389 77 2405 111
rect 2339 61 2405 77
rect 2357 39 2387 61
rect 2357 -183 2387 -161
rect 2339 -199 2405 -183
rect 2339 -233 2355 -199
rect 2389 -233 2405 -199
rect 2339 -249 2405 -233
rect 2708 76 2774 92
rect 2708 42 2724 76
rect 2758 42 2774 76
rect 2708 26 2774 42
rect 2726 -5 2756 26
rect 2726 -232 2756 -205
rect -10 -404 56 -388
rect -10 -438 6 -404
rect 40 -438 56 -404
rect -10 -454 56 -438
rect 3077 23 3143 39
rect 3077 -11 3093 23
rect 3127 -11 3143 23
rect 3077 -27 3143 -11
rect 3095 -58 3125 -27
rect 3095 -285 3125 -258
rect 8 -476 38 -454
rect 8 -902 38 -876
rect 3446 -30 3512 -14
rect 3446 -64 3462 -30
rect 3496 -64 3512 -30
rect 3446 -80 3512 -64
rect 3464 -111 3494 -80
rect 3464 -338 3494 -311
rect 3815 -101 3881 -85
rect 3815 -135 3831 -101
rect 3865 -135 3881 -101
rect 3815 -151 3881 -135
rect 3833 -173 3863 -151
rect 3833 -395 3863 -373
rect 3815 -411 3881 -395
rect 3815 -445 3831 -411
rect 3865 -445 3881 -411
rect 3815 -461 3881 -445
rect 4184 -154 4250 -138
rect 4184 -188 4200 -154
rect 4234 -188 4250 -154
rect 4184 -204 4250 -188
rect 4202 -226 4232 -204
rect 4202 -448 4232 -426
rect 4184 -464 4250 -448
rect 4184 -498 4200 -464
rect 4234 -498 4250 -464
rect 4184 -514 4250 -498
rect 4553 -207 4619 -191
rect 4553 -241 4569 -207
rect 4603 -241 4619 -207
rect 4553 -257 4619 -241
rect 4571 -279 4601 -257
rect 4571 -501 4601 -479
rect 4553 -517 4619 -501
rect 4553 -551 4569 -517
rect 4603 -551 4619 -517
rect 4553 -567 4619 -551
rect 4922 -242 4988 -226
rect 4922 -276 4938 -242
rect 4972 -276 4988 -242
rect 4922 -292 4988 -276
rect 4940 -323 4970 -292
rect 4940 -550 4970 -523
rect 5291 -295 5357 -279
rect 5291 -329 5307 -295
rect 5341 -329 5357 -295
rect 5291 -345 5357 -329
rect 5309 -376 5339 -345
rect 5309 -603 5339 -576
rect 5660 -348 5726 -332
rect 5660 -382 5676 -348
rect 5710 -382 5726 -348
rect 5660 -398 5726 -382
rect 5678 -429 5708 -398
rect 5678 -656 5708 -629
rect 6029 -419 6095 -403
rect 6029 -453 6045 -419
rect 6079 -453 6095 -419
rect 6029 -469 6095 -453
rect 6047 -491 6077 -469
rect 6047 -713 6077 -691
rect 6029 -729 6095 -713
rect 6029 -763 6045 -729
rect 6079 -763 6095 -729
rect 6029 -779 6095 -763
rect 6398 -472 6464 -456
rect 6398 -506 6414 -472
rect 6448 -506 6464 -472
rect 6398 -522 6464 -506
rect 6416 -544 6446 -522
rect 6416 -766 6446 -744
rect 6398 -782 6464 -766
rect 6398 -816 6414 -782
rect 6448 -816 6464 -782
rect 6398 -832 6464 -816
rect 6767 -525 6833 -509
rect 6767 -559 6783 -525
rect 6817 -559 6833 -525
rect 6767 -575 6833 -559
rect 6785 -597 6815 -575
rect 6785 -819 6815 -797
rect 6767 -835 6833 -819
rect 6767 -869 6783 -835
rect 6817 -869 6833 -835
rect 6767 -885 6833 -869
rect 7136 -560 7202 -544
rect 7136 -594 7152 -560
rect 7186 -594 7202 -560
rect 7136 -610 7202 -594
rect 7154 -641 7184 -610
rect 7154 -868 7184 -841
rect 7505 -613 7571 -597
rect 7505 -647 7521 -613
rect 7555 -647 7571 -613
rect 7505 -663 7571 -647
rect 7523 -694 7553 -663
rect 7523 -921 7553 -894
rect 7874 -666 7940 -650
rect 7874 -700 7890 -666
rect 7924 -700 7940 -666
rect 7874 -716 7940 -700
rect 7892 -747 7922 -716
rect 7892 -974 7922 -947
rect 8243 -737 8309 -721
rect 8243 -771 8259 -737
rect 8293 -771 8309 -737
rect 8243 -787 8309 -771
rect 8261 -809 8291 -787
rect 8261 -1031 8291 -1009
rect 8243 -1047 8309 -1031
rect 8243 -1081 8259 -1047
rect 8293 -1081 8309 -1047
rect 8243 -1097 8309 -1081
<< polycont >>
rect -540 644 -506 678
rect 504 416 538 450
rect -418 -80 -384 -46
rect 998 408 1032 442
rect 998 98 1032 132
rect 1986 130 2020 164
rect 1986 -180 2020 -146
rect 2355 77 2389 111
rect 2355 -233 2389 -199
rect 2724 42 2758 76
rect 6 -438 40 -404
rect 3093 -11 3127 23
rect 3462 -64 3496 -30
rect 3831 -135 3865 -101
rect 3831 -445 3865 -411
rect 4200 -188 4234 -154
rect 4200 -498 4234 -464
rect 4569 -241 4603 -207
rect 4569 -551 4603 -517
rect 4938 -276 4972 -242
rect 5307 -329 5341 -295
rect 5676 -382 5710 -348
rect 6045 -453 6079 -419
rect 6045 -763 6079 -729
rect 6414 -506 6448 -472
rect 6414 -816 6448 -782
rect 6783 -559 6817 -525
rect 6783 -869 6817 -835
rect 7152 -594 7186 -560
rect 7521 -647 7555 -613
rect 7890 -700 7924 -666
rect 8259 -771 8293 -737
rect 8259 -1081 8293 -1047
<< locali >>
rect -698 746 -602 780
rect -444 746 -348 780
rect -698 684 -664 746
rect -382 684 -348 746
rect -584 644 -540 678
rect -506 644 -490 678
rect -584 585 -550 644
rect -584 393 -550 409
rect -496 585 -462 601
rect -496 393 -462 409
rect -698 248 -664 310
rect -382 248 -348 310
rect -698 214 -602 248
rect -444 214 -348 248
rect 346 518 442 552
rect 600 518 696 552
rect 346 456 380 518
rect 662 456 696 518
rect 488 416 504 450
rect 538 416 554 450
rect 460 357 494 373
rect 460 165 494 181
rect 548 357 582 373
rect 548 165 582 181
rect -576 22 -480 56
rect -322 22 -226 56
rect -576 -40 -542 22
rect -260 -40 -226 22
rect 346 20 380 82
rect 662 20 696 82
rect 346 -14 442 20
rect 600 -14 696 20
rect 840 510 936 544
rect 1094 510 1190 544
rect 840 448 874 510
rect 1156 448 1190 510
rect 982 408 998 442
rect 1032 408 1048 442
rect 954 358 988 374
rect 954 166 988 182
rect 1042 358 1076 374
rect 1042 166 1076 182
rect 982 98 998 132
rect 1032 98 1048 132
rect 840 30 874 92
rect 1156 30 1190 92
rect 840 -4 936 30
rect 1094 -4 1190 30
rect 1828 232 1924 266
rect 2082 232 2178 266
rect 1828 170 1862 232
rect -434 -80 -418 -46
rect -384 -80 -368 -46
rect -462 -130 -428 -114
rect -462 -522 -428 -506
rect -374 -130 -340 -114
rect -374 -522 -340 -506
rect -576 -658 -542 -596
rect 2144 170 2178 232
rect 1970 130 1986 164
rect 2020 130 2036 164
rect 1942 80 1976 96
rect 1942 -112 1976 -96
rect 2030 80 2064 96
rect 2030 -112 2064 -96
rect 1970 -180 1986 -146
rect 2020 -180 2036 -146
rect 1828 -248 1862 -186
rect 2144 -248 2178 -186
rect 1828 -282 1924 -248
rect 2082 -282 2178 -248
rect 2197 179 2293 213
rect 2451 179 2547 213
rect 2197 117 2231 179
rect 2513 117 2547 179
rect 2339 77 2355 111
rect 2389 77 2405 111
rect 2311 27 2345 43
rect 2311 -165 2345 -149
rect 2399 27 2433 43
rect 2399 -165 2433 -149
rect 2339 -233 2355 -199
rect 2389 -233 2405 -199
rect 2197 -301 2231 -239
rect 2513 -301 2547 -239
rect -260 -658 -226 -596
rect -576 -692 -480 -658
rect -322 -692 -226 -658
rect -152 -336 -56 -302
rect 102 -336 198 -302
rect 2197 -335 2293 -301
rect 2451 -335 2547 -301
rect 2566 144 2662 178
rect 2820 144 2916 178
rect 2566 82 2600 144
rect 2882 82 2916 144
rect 2708 42 2724 76
rect 2758 42 2774 76
rect 2680 -17 2714 -1
rect 2680 -209 2714 -193
rect 2768 -17 2802 -1
rect 2768 -209 2802 -193
rect -152 -398 -118 -336
rect 164 -398 198 -336
rect 2566 -354 2600 -292
rect 2882 -354 2916 -292
rect 2566 -388 2662 -354
rect 2820 -388 2916 -354
rect 2935 91 3031 125
rect 3189 91 3285 125
rect 2935 29 2969 91
rect 3251 29 3285 91
rect 3077 -11 3093 23
rect 3127 -11 3143 23
rect 3049 -70 3083 -54
rect 3049 -262 3083 -246
rect 3137 -70 3171 -54
rect 3137 -262 3171 -246
rect -38 -438 6 -404
rect 40 -438 56 -404
rect -38 -472 -2 -438
rect -38 -488 -4 -472
rect -38 -880 -4 -864
rect 50 -488 84 -472
rect 50 -880 84 -864
rect -152 -1016 -118 -954
rect 2935 -407 2969 -345
rect 3251 -407 3285 -345
rect 2935 -441 3031 -407
rect 3189 -441 3285 -407
rect 3304 38 3400 72
rect 3558 38 3654 72
rect 3304 -24 3338 38
rect 3620 -24 3654 38
rect 3446 -64 3462 -30
rect 3496 -64 3512 -30
rect 3418 -123 3452 -107
rect 3418 -315 3452 -299
rect 3506 -123 3540 -107
rect 3506 -315 3540 -299
rect 3304 -460 3338 -398
rect 3620 -460 3654 -398
rect 3304 -494 3400 -460
rect 3558 -494 3654 -460
rect 3673 -33 3769 1
rect 3927 -33 4023 1
rect 3673 -95 3707 -33
rect 3989 -95 4023 -33
rect 3815 -135 3831 -101
rect 3865 -135 3881 -101
rect 3787 -185 3821 -169
rect 3787 -377 3821 -361
rect 3875 -185 3909 -169
rect 3875 -377 3909 -361
rect 3815 -445 3831 -411
rect 3865 -445 3881 -411
rect 3673 -513 3707 -451
rect 3989 -513 4023 -451
rect 3673 -547 3769 -513
rect 3927 -547 4023 -513
rect 4042 -86 4138 -52
rect 4296 -86 4392 -52
rect 4042 -148 4076 -86
rect 4358 -148 4392 -86
rect 4184 -188 4200 -154
rect 4234 -188 4250 -154
rect 4156 -238 4190 -222
rect 4156 -430 4190 -414
rect 4244 -238 4278 -222
rect 4244 -430 4278 -414
rect 4184 -498 4200 -464
rect 4234 -498 4250 -464
rect 4042 -566 4076 -504
rect 4358 -566 4392 -504
rect 4042 -600 4138 -566
rect 4296 -600 4392 -566
rect 4411 -139 4507 -105
rect 4665 -139 4761 -105
rect 4411 -201 4445 -139
rect 4727 -201 4761 -139
rect 4553 -241 4569 -207
rect 4603 -241 4619 -207
rect 4525 -291 4559 -275
rect 4525 -483 4559 -467
rect 4613 -291 4647 -275
rect 4613 -483 4647 -467
rect 4553 -551 4569 -517
rect 4603 -551 4619 -517
rect 4411 -619 4445 -557
rect 4727 -619 4761 -557
rect 4411 -653 4507 -619
rect 4665 -653 4761 -619
rect 4780 -174 4876 -140
rect 5034 -174 5130 -140
rect 4780 -236 4814 -174
rect 5096 -236 5130 -174
rect 4922 -276 4938 -242
rect 4972 -276 4988 -242
rect 4894 -335 4928 -319
rect 4894 -527 4928 -511
rect 4982 -335 5016 -319
rect 4982 -527 5016 -511
rect 4780 -672 4814 -610
rect 5096 -672 5130 -610
rect 4780 -706 4876 -672
rect 5034 -706 5130 -672
rect 5149 -227 5245 -193
rect 5403 -227 5499 -193
rect 5149 -289 5183 -227
rect 5465 -289 5499 -227
rect 5291 -329 5307 -295
rect 5341 -329 5357 -295
rect 5263 -388 5297 -372
rect 5263 -580 5297 -564
rect 5351 -388 5385 -372
rect 5351 -580 5385 -564
rect 5149 -725 5183 -663
rect 5465 -725 5499 -663
rect 5149 -759 5245 -725
rect 5403 -759 5499 -725
rect 5518 -280 5614 -246
rect 5772 -280 5868 -246
rect 5518 -342 5552 -280
rect 5834 -342 5868 -280
rect 5660 -382 5676 -348
rect 5710 -382 5726 -348
rect 5632 -441 5666 -425
rect 5632 -633 5666 -617
rect 5720 -441 5754 -425
rect 5720 -633 5754 -617
rect 5518 -778 5552 -716
rect 5834 -778 5868 -716
rect 5518 -812 5614 -778
rect 5772 -812 5868 -778
rect 5887 -351 5983 -317
rect 6141 -351 6237 -317
rect 5887 -413 5921 -351
rect 6203 -413 6237 -351
rect 6029 -453 6045 -419
rect 6079 -453 6095 -419
rect 6001 -503 6035 -487
rect 6001 -695 6035 -679
rect 6089 -503 6123 -487
rect 6089 -695 6123 -679
rect 6029 -763 6045 -729
rect 6079 -763 6095 -729
rect 5887 -831 5921 -769
rect 6203 -831 6237 -769
rect 5887 -865 5983 -831
rect 6141 -865 6237 -831
rect 6256 -404 6352 -370
rect 6510 -404 6606 -370
rect 6256 -466 6290 -404
rect 6572 -466 6606 -404
rect 6398 -506 6414 -472
rect 6448 -506 6464 -472
rect 6370 -556 6404 -540
rect 6370 -748 6404 -732
rect 6458 -556 6492 -540
rect 6458 -748 6492 -732
rect 6398 -816 6414 -782
rect 6448 -816 6464 -782
rect 6256 -884 6290 -822
rect 6572 -884 6606 -822
rect 6256 -918 6352 -884
rect 6510 -918 6606 -884
rect 6625 -457 6721 -423
rect 6879 -457 6975 -423
rect 6625 -519 6659 -457
rect 6941 -519 6975 -457
rect 6767 -559 6783 -525
rect 6817 -559 6833 -525
rect 6739 -609 6773 -593
rect 6739 -801 6773 -785
rect 6827 -609 6861 -593
rect 6827 -801 6861 -785
rect 6767 -869 6783 -835
rect 6817 -869 6833 -835
rect 164 -1016 198 -954
rect 6625 -937 6659 -875
rect 6941 -937 6975 -875
rect 6625 -971 6721 -937
rect 6879 -971 6975 -937
rect 6994 -492 7090 -458
rect 7248 -492 7344 -458
rect 6994 -554 7028 -492
rect 7310 -554 7344 -492
rect 7136 -594 7152 -560
rect 7186 -594 7202 -560
rect 7108 -653 7142 -637
rect 7108 -845 7142 -829
rect 7196 -653 7230 -637
rect 7196 -845 7230 -829
rect -152 -1050 -56 -1016
rect 102 -1050 198 -1016
rect 6994 -990 7028 -928
rect 7310 -990 7344 -928
rect 6994 -1024 7090 -990
rect 7248 -1024 7344 -990
rect 7363 -545 7459 -511
rect 7617 -545 7713 -511
rect 7363 -607 7397 -545
rect 7679 -607 7713 -545
rect 7505 -647 7521 -613
rect 7555 -647 7571 -613
rect 7477 -706 7511 -690
rect 7477 -898 7511 -882
rect 7565 -706 7599 -690
rect 7565 -898 7599 -882
rect 7363 -1043 7397 -981
rect 7679 -1043 7713 -981
rect 7363 -1077 7459 -1043
rect 7617 -1077 7713 -1043
rect 7732 -598 7828 -564
rect 7986 -598 8082 -564
rect 7732 -660 7766 -598
rect 8048 -660 8082 -598
rect 7874 -700 7890 -666
rect 7924 -700 7940 -666
rect 7846 -759 7880 -743
rect 7846 -951 7880 -935
rect 7934 -759 7968 -743
rect 7934 -951 7968 -935
rect 7732 -1096 7766 -1034
rect 8048 -1096 8082 -1034
rect 7732 -1130 7828 -1096
rect 7986 -1130 8082 -1096
rect 8101 -669 8197 -635
rect 8355 -669 8451 -635
rect 8101 -731 8135 -669
rect 8417 -731 8451 -669
rect 8243 -771 8259 -737
rect 8293 -771 8309 -737
rect 8215 -821 8249 -805
rect 8215 -1013 8249 -997
rect 8303 -821 8337 -805
rect 8303 -1013 8337 -997
rect 8243 -1081 8259 -1047
rect 8293 -1081 8309 -1047
rect 8101 -1149 8135 -1087
rect 8417 -1149 8451 -1087
rect 8101 -1183 8197 -1149
rect 8355 -1183 8451 -1149
<< viali >>
rect -540 644 -506 678
rect -584 409 -550 585
rect -496 409 -462 585
rect 504 416 538 450
rect 460 181 494 357
rect 548 181 582 357
rect 998 408 1032 442
rect 954 182 988 358
rect 1042 182 1076 358
rect 998 98 1032 132
rect -418 -80 -384 -46
rect -462 -506 -428 -130
rect -374 -506 -340 -130
rect 1986 130 2020 164
rect 1942 -96 1976 80
rect 2030 -96 2064 80
rect 1986 -180 2020 -146
rect 2355 77 2389 111
rect 2311 -149 2345 27
rect 2399 -149 2433 27
rect 2355 -233 2389 -199
rect 2724 42 2758 76
rect 2680 -193 2714 -17
rect 2768 -193 2802 -17
rect 3093 -11 3127 23
rect 3049 -246 3083 -70
rect 3137 -246 3171 -70
rect 6 -438 40 -404
rect -38 -864 -4 -488
rect 50 -864 84 -488
rect 3462 -64 3496 -30
rect 3418 -299 3452 -123
rect 3506 -299 3540 -123
rect 3831 -135 3865 -101
rect 3787 -361 3821 -185
rect 3875 -361 3909 -185
rect 3831 -445 3865 -411
rect 4200 -188 4234 -154
rect 4156 -414 4190 -238
rect 4244 -414 4278 -238
rect 4200 -498 4234 -464
rect 4569 -241 4603 -207
rect 4525 -467 4559 -291
rect 4613 -467 4647 -291
rect 4569 -551 4603 -517
rect 4938 -276 4972 -242
rect 4894 -511 4928 -335
rect 4982 -511 5016 -335
rect 5307 -329 5341 -295
rect 5263 -564 5297 -388
rect 5351 -564 5385 -388
rect 5676 -382 5710 -348
rect 5632 -617 5666 -441
rect 5720 -617 5754 -441
rect 6045 -453 6079 -419
rect 6001 -679 6035 -503
rect 6089 -679 6123 -503
rect 6045 -763 6079 -729
rect 6414 -506 6448 -472
rect 6370 -732 6404 -556
rect 6458 -732 6492 -556
rect 6414 -816 6448 -782
rect 6783 -559 6817 -525
rect 6739 -785 6773 -609
rect 6827 -785 6861 -609
rect 6783 -869 6817 -835
rect 7152 -594 7186 -560
rect 7108 -829 7142 -653
rect 7196 -829 7230 -653
rect 7521 -647 7555 -613
rect 7477 -882 7511 -706
rect 7565 -882 7599 -706
rect 7890 -700 7924 -666
rect 7846 -935 7880 -759
rect 7934 -935 7968 -759
rect 8259 -771 8293 -737
rect 8215 -997 8249 -821
rect 8303 -997 8337 -821
rect 8259 -1081 8293 -1047
<< metal1 >>
rect -856 726 -212 802
rect -552 678 -492 690
rect -552 644 -540 678
rect -506 644 -492 678
rect -552 634 -492 644
rect -496 597 -60 604
rect -590 585 -544 597
rect -590 409 -584 585
rect -550 409 -544 585
rect -590 397 -544 409
rect -502 585 -60 597
rect -502 409 -496 585
rect -462 554 -60 585
rect -462 409 -456 554
rect 542 456 994 468
rect 492 450 994 456
rect 492 416 504 450
rect 538 448 994 450
rect 538 442 1044 448
rect 538 416 998 442
rect 492 410 998 416
rect -502 397 -456 409
rect 542 408 998 410
rect 1032 408 1044 442
rect 542 402 1044 408
rect -584 -118 -550 397
rect 454 357 500 369
rect 454 181 460 357
rect 494 181 500 357
rect 454 169 500 181
rect 542 357 588 369
rect 542 181 548 357
rect 582 181 588 357
rect 542 169 588 181
rect 948 358 994 370
rect 948 182 954 358
rect 988 182 994 358
rect 948 170 994 182
rect 1036 358 1082 370
rect 1036 182 1042 358
rect 1076 182 1082 358
rect 1036 170 1082 182
rect 1974 164 2032 170
rect 986 132 1044 138
rect 986 98 998 132
rect 1032 98 1044 132
rect 1974 130 1986 164
rect 2020 130 2032 164
rect 1974 124 2032 130
rect 986 92 1044 98
rect 2343 111 2401 117
rect 1936 80 1982 92
rect -346 -34 -98 -32
rect -404 -40 -98 -34
rect -430 -46 -98 -40
rect -430 -80 -418 -46
rect -384 -80 -98 -46
rect -430 -86 -98 -80
rect -346 -88 -98 -86
rect 1936 -96 1942 80
rect 1976 -96 1982 80
rect 1936 -108 1982 -96
rect 2024 80 2070 92
rect 2024 -96 2030 80
rect 2064 -96 2070 80
rect 2343 77 2355 111
rect 2389 77 2401 111
rect 2343 71 2401 77
rect 2712 76 2770 82
rect 2712 42 2724 76
rect 2758 42 2770 76
rect 2024 -108 2070 -96
rect 2305 27 2351 39
rect -584 -130 -422 -118
rect -584 -162 -462 -130
rect -468 -506 -462 -162
rect -428 -506 -422 -130
rect -468 -518 -422 -506
rect -380 -130 -334 -118
rect -380 -506 -374 -130
rect -340 -474 -334 -130
rect 1974 -146 2032 -140
rect 1974 -180 1986 -146
rect 2020 -180 2032 -146
rect 2305 -149 2311 27
rect 2345 -149 2351 27
rect 2305 -161 2351 -149
rect 2393 27 2439 39
rect 2712 36 2770 42
rect 2393 -149 2399 27
rect 2433 -149 2439 27
rect 3081 23 3139 29
rect 2393 -161 2439 -149
rect 2674 -17 2720 -5
rect 1974 -186 2032 -180
rect 2674 -193 2680 -17
rect 2714 -193 2720 -17
rect 2343 -199 2401 -193
rect 2343 -233 2355 -199
rect 2389 -233 2401 -199
rect 2674 -205 2720 -193
rect 2762 -17 2808 -5
rect 3081 -11 3093 23
rect 3127 -11 3139 23
rect 3081 -17 3139 -11
rect 2762 -193 2768 -17
rect 2802 -193 2808 -17
rect 3450 -30 3508 -24
rect 2762 -205 2808 -193
rect 3043 -70 3089 -58
rect 2343 -239 2401 -233
rect 3043 -246 3049 -70
rect 3083 -246 3089 -70
rect 3043 -258 3089 -246
rect 3131 -70 3177 -58
rect 3450 -64 3462 -30
rect 3496 -64 3508 -30
rect 3450 -70 3508 -64
rect 3131 -246 3137 -70
rect 3171 -246 3177 -70
rect 3819 -101 3877 -95
rect 3131 -258 3177 -246
rect 3412 -123 3458 -111
rect 3412 -299 3418 -123
rect 3452 -299 3458 -123
rect 3412 -311 3458 -299
rect 3500 -123 3546 -111
rect 3500 -299 3506 -123
rect 3540 -299 3546 -123
rect 3819 -135 3831 -101
rect 3865 -135 3877 -101
rect 3819 -141 3877 -135
rect 4188 -154 4246 -148
rect 3500 -311 3546 -299
rect 3781 -185 3827 -173
rect 3781 -361 3787 -185
rect 3821 -361 3827 -185
rect 3781 -373 3827 -361
rect 3869 -185 3915 -173
rect 3869 -361 3875 -185
rect 3909 -361 3915 -185
rect 4188 -188 4200 -154
rect 4234 -188 4246 -154
rect 4188 -194 4246 -188
rect 4557 -207 4615 -201
rect 3869 -373 3915 -361
rect 4150 -238 4196 -226
rect -8 -404 54 -392
rect -8 -438 6 -404
rect 40 -438 54 -404
rect -8 -446 54 -438
rect 3819 -411 3877 -405
rect 3819 -445 3831 -411
rect 3865 -445 3877 -411
rect 4150 -414 4156 -238
rect 4190 -414 4196 -238
rect 4150 -426 4196 -414
rect 4238 -238 4284 -226
rect 4238 -414 4244 -238
rect 4278 -414 4284 -238
rect 4557 -241 4569 -207
rect 4603 -241 4615 -207
rect 4557 -247 4615 -241
rect 4926 -242 4984 -236
rect 4926 -276 4938 -242
rect 4972 -276 4984 -242
rect 4238 -426 4284 -414
rect 4519 -291 4565 -279
rect 3819 -451 3877 -445
rect 4188 -464 4246 -458
rect -340 -488 4 -474
rect -340 -506 -38 -488
rect -380 -554 -38 -506
rect -44 -864 -38 -554
rect -4 -554 4 -488
rect 44 -488 90 -476
rect -4 -864 2 -554
rect -44 -876 2 -864
rect 44 -864 50 -488
rect 84 -864 90 -488
rect 4188 -498 4200 -464
rect 4234 -498 4246 -464
rect 4519 -467 4525 -291
rect 4559 -467 4565 -291
rect 4519 -479 4565 -467
rect 4607 -291 4653 -279
rect 4926 -282 4984 -276
rect 4607 -467 4613 -291
rect 4647 -467 4653 -291
rect 5295 -295 5353 -289
rect 4607 -479 4653 -467
rect 4888 -335 4934 -323
rect 4188 -504 4246 -498
rect 4888 -511 4894 -335
rect 4928 -511 4934 -335
rect 4557 -517 4615 -511
rect 4557 -551 4569 -517
rect 4603 -551 4615 -517
rect 4888 -523 4934 -511
rect 4976 -335 5022 -323
rect 5295 -329 5307 -295
rect 5341 -329 5353 -295
rect 5295 -335 5353 -329
rect 4976 -511 4982 -335
rect 5016 -511 5022 -335
rect 5664 -348 5722 -342
rect 4976 -523 5022 -511
rect 5257 -388 5303 -376
rect 4557 -557 4615 -551
rect 5257 -564 5263 -388
rect 5297 -564 5303 -388
rect 5257 -576 5303 -564
rect 5345 -388 5391 -376
rect 5664 -382 5676 -348
rect 5710 -382 5722 -348
rect 5664 -388 5722 -382
rect 5345 -564 5351 -388
rect 5385 -564 5391 -388
rect 6033 -419 6091 -413
rect 5345 -576 5391 -564
rect 5626 -441 5672 -429
rect 5626 -617 5632 -441
rect 5666 -617 5672 -441
rect 5626 -629 5672 -617
rect 5714 -441 5760 -429
rect 5714 -617 5720 -441
rect 5754 -617 5760 -441
rect 6033 -453 6045 -419
rect 6079 -453 6091 -419
rect 6033 -459 6091 -453
rect 6402 -472 6460 -466
rect 5714 -629 5760 -617
rect 5995 -503 6041 -491
rect 5995 -679 6001 -503
rect 6035 -679 6041 -503
rect 5995 -691 6041 -679
rect 6083 -503 6129 -491
rect 6083 -679 6089 -503
rect 6123 -679 6129 -503
rect 6402 -506 6414 -472
rect 6448 -506 6460 -472
rect 6402 -512 6460 -506
rect 6771 -525 6829 -519
rect 6083 -691 6129 -679
rect 6364 -556 6410 -544
rect 6033 -729 6091 -723
rect 6033 -763 6045 -729
rect 6079 -763 6091 -729
rect 6364 -732 6370 -556
rect 6404 -732 6410 -556
rect 6364 -744 6410 -732
rect 6452 -556 6498 -544
rect 6452 -732 6458 -556
rect 6492 -732 6498 -556
rect 6771 -559 6783 -525
rect 6817 -559 6829 -525
rect 6771 -565 6829 -559
rect 7140 -560 7198 -554
rect 7140 -594 7152 -560
rect 7186 -594 7198 -560
rect 6452 -744 6498 -732
rect 6733 -609 6779 -597
rect 6033 -769 6091 -763
rect 6402 -782 6460 -776
rect 6402 -816 6414 -782
rect 6448 -816 6460 -782
rect 6733 -785 6739 -609
rect 6773 -785 6779 -609
rect 6733 -797 6779 -785
rect 6821 -609 6867 -597
rect 7140 -600 7198 -594
rect 6821 -785 6827 -609
rect 6861 -785 6867 -609
rect 7509 -613 7567 -607
rect 6821 -797 6867 -785
rect 7102 -653 7148 -641
rect 6402 -822 6460 -816
rect 7102 -829 7108 -653
rect 7142 -829 7148 -653
rect 44 -876 90 -864
rect 6771 -835 6829 -829
rect 6771 -869 6783 -835
rect 6817 -869 6829 -835
rect 7102 -841 7148 -829
rect 7190 -653 7236 -641
rect 7509 -647 7521 -613
rect 7555 -647 7567 -613
rect 7509 -653 7567 -647
rect 7190 -829 7196 -653
rect 7230 -829 7236 -653
rect 7878 -666 7936 -660
rect 7190 -841 7236 -829
rect 7471 -706 7517 -694
rect 6771 -875 6829 -869
rect 7471 -882 7477 -706
rect 7511 -882 7517 -706
rect 7471 -894 7517 -882
rect 7559 -706 7605 -694
rect 7878 -700 7890 -666
rect 7924 -700 7936 -666
rect 7878 -706 7936 -700
rect 7559 -882 7565 -706
rect 7599 -882 7605 -706
rect 8247 -737 8305 -731
rect 7559 -894 7605 -882
rect 7840 -759 7886 -747
rect 7840 -935 7846 -759
rect 7880 -935 7886 -759
rect 7840 -947 7886 -935
rect 7928 -759 7974 -747
rect 7928 -935 7934 -759
rect 7968 -935 7974 -759
rect 8247 -771 8259 -737
rect 8293 -771 8305 -737
rect 8247 -777 8305 -771
rect 7928 -947 7974 -935
rect 8209 -821 8255 -809
rect 8209 -997 8215 -821
rect 8249 -997 8255 -821
rect 8209 -1009 8255 -997
rect 8297 -821 8343 -809
rect 8297 -997 8303 -821
rect 8337 -997 8343 -821
rect 8297 -1009 8343 -997
rect 8247 -1047 8305 -1041
rect 8247 -1081 8259 -1047
rect 8293 -1081 8305 -1047
rect 8247 -1087 8305 -1081
<< labels >>
rlabel psubdiffcont 23 -1033 23 -1033 0 XM2.B
rlabel ndiffc -21 -676 -21 -676 0 XM2.D
rlabel ndiffc 67 -676 67 -676 0 XM2.S
rlabel polycont 23 -421 23 -421 0 XM2.G
rlabel psubdiffcont -401 -675 -401 -675 0 XM1.B
rlabel ndiffc -445 -318 -445 -318 0 XM1.D
rlabel ndiffc -357 -318 -357 -318 0 XM1.S
rlabel polycont -401 -63 -401 -63 0 XM1.G
rlabel psubdiffcont 2003 -265 2003 -265 0 XM11.B
rlabel ndiffc 1959 -8 1959 -8 0 XM11.D
rlabel ndiffc 2047 -8 2047 -8 0 XM11.S
rlabel polycont 2003 147 2003 147 0 XM11.G
rlabel psubdiffcont 2372 -318 2372 -318 0 XM12.B
rlabel ndiffc 2328 -61 2328 -61 0 XM12.D
rlabel ndiffc 2416 -61 2416 -61 0 XM12.S
rlabel polycont 2372 94 2372 94 0 XM12.G
rlabel nsubdiffcont 2741 -371 2741 -371 0 XM13.B
rlabel pdiffc 2697 -105 2697 -105 0 XM13.D
rlabel pdiffc 2785 -105 2785 -105 0 XM13.S
rlabel polycont 2741 59 2741 59 0 XM13.G
rlabel nsubdiffcont 3110 -424 3110 -424 0 XM14.B
rlabel pdiffc 3066 -158 3066 -158 0 XM14.D
rlabel pdiffc 3154 -158 3154 -158 0 XM14.S
rlabel polycont 3110 6 3110 6 0 XM14.G
rlabel nsubdiffcont 3479 -477 3479 -477 0 XM19.B
rlabel pdiffc 3435 -211 3435 -211 0 XM19.D
rlabel pdiffc 3523 -211 3523 -211 0 XM19.S
rlabel polycont 3479 -47 3479 -47 0 XM19.G
rlabel psubdiffcont 3848 -530 3848 -530 0 XM20.B
rlabel ndiffc 3804 -273 3804 -273 0 XM20.D
rlabel ndiffc 3892 -273 3892 -273 0 XM20.S
rlabel polycont 3848 -118 3848 -118 0 XM20.G
rlabel psubdiffcont 4217 -583 4217 -583 0 XM21.B
rlabel ndiffc 4173 -326 4173 -326 0 XM21.D
rlabel ndiffc 4261 -326 4261 -326 0 XM21.S
rlabel polycont 4217 -171 4217 -171 0 XM21.G
rlabel psubdiffcont 4586 -636 4586 -636 0 XM22.B
rlabel ndiffc 4542 -379 4542 -379 0 XM22.D
rlabel ndiffc 4630 -379 4630 -379 0 XM22.S
rlabel polycont 4586 -224 4586 -224 0 XM22.G
rlabel nsubdiffcont 4955 -689 4955 -689 0 XM23.B
rlabel pdiffc 4911 -423 4911 -423 0 XM23.D
rlabel pdiffc 4999 -423 4999 -423 0 XM23.S
rlabel polycont 4955 -259 4955 -259 0 XM23.G
rlabel nsubdiffcont 5324 -742 5324 -742 0 XM24.B
rlabel pdiffc 5280 -476 5280 -476 0 XM24.D
rlabel pdiffc 5368 -476 5368 -476 0 XM24.S
rlabel polycont 5324 -312 5324 -312 0 XM24.G
rlabel nsubdiffcont 5693 -795 5693 -795 0 XM25.B
rlabel pdiffc 5649 -529 5649 -529 0 XM25.D
rlabel pdiffc 5737 -529 5737 -529 0 XM25.S
rlabel polycont 5693 -365 5693 -365 0 XM25.G
rlabel psubdiffcont 6062 -848 6062 -848 0 XM26.B
rlabel ndiffc 6018 -591 6018 -591 0 XM26.D
rlabel ndiffc 6106 -591 6106 -591 0 XM26.S
rlabel polycont 6062 -436 6062 -436 0 XM26.G
rlabel psubdiffcont 6431 -901 6431 -901 0 XM27.B
rlabel ndiffc 6387 -644 6387 -644 0 XM27.D
rlabel ndiffc 6475 -644 6475 -644 0 XM27.S
rlabel polycont 6431 -489 6431 -489 0 XM27.G
rlabel psubdiffcont 6800 -954 6800 -954 0 XM28.B
rlabel ndiffc 6756 -697 6756 -697 0 XM28.D
rlabel ndiffc 6844 -697 6844 -697 0 XM28.S
rlabel polycont 6800 -542 6800 -542 0 XM28.G
rlabel nsubdiffcont 7169 -1007 7169 -1007 0 XM29.B
rlabel pdiffc 7125 -741 7125 -741 0 XM29.D
rlabel pdiffc 7213 -741 7213 -741 0 XM29.S
rlabel polycont 7169 -577 7169 -577 0 XM29.G
rlabel nsubdiffcont 7538 -1060 7538 -1060 0 XM30.B
rlabel pdiffc 7494 -794 7494 -794 0 XM30.D
rlabel pdiffc 7582 -794 7582 -794 0 XM30.S
rlabel polycont 7538 -630 7538 -630 0 XM30.G
rlabel nsubdiffcont 7907 -1113 7907 -1113 0 XM31.B
rlabel pdiffc 7863 -847 7863 -847 0 XM31.D
rlabel pdiffc 7951 -847 7951 -847 0 XM31.S
rlabel polycont 7907 -683 7907 -683 0 XM31.G
rlabel psubdiffcont 8276 -1166 8276 -1166 0 XM32.B
rlabel ndiffc 8232 -909 8232 -909 0 XM32.D
rlabel ndiffc 8320 -909 8320 -909 0 XM32.S
rlabel polycont 8276 -754 8276 -754 0 XM32.G
rlabel nsubdiffcont -523 231 -523 231 0 XM3.B
rlabel pdiffc -567 497 -567 497 0 XM3.D
rlabel pdiffc -479 497 -479 497 0 XM3.S
rlabel polycont -523 661 -523 661 0 XM3.G
rlabel psubdiffcont 1015 13 1015 13 0 XM4.B
rlabel ndiffc 971 270 971 270 0 XM4.D
rlabel ndiffc 1059 270 1059 270 0 XM4.S
rlabel polycont 1015 425 1015 425 0 XM4.G
rlabel nsubdiffcont 521 3 521 3 0 XM5.B
rlabel pdiffc 477 269 477 269 0 XM5.D
rlabel pdiffc 565 269 565 269 0 XM5.S
rlabel polycont 521 433 521 433 0 XM5.G
<< end >>
