magic
tech sky130A
magscale 1 2
timestamp 1745430941
<< locali >>
rect 5926 1510 6120 1518
rect 5124 1506 6120 1510
rect -668 1452 6120 1506
rect -668 1418 -493 1452
rect -387 1418 6120 1452
rect -668 1336 6120 1418
rect -668 1288 268 1336
rect -668 740 -480 1288
rect -100 1274 268 1288
rect -100 792 266 1274
rect 592 792 958 1336
rect 1684 794 2042 1336
rect 2364 794 2718 1336
rect 1684 792 2718 794
rect 3444 814 3794 1336
rect 4124 814 4468 1336
rect 5204 814 5566 1336
rect 5592 1332 6120 1336
rect 5894 814 6120 1332
rect 3444 792 6120 814
rect -100 740 6120 792
rect -668 536 6120 740
rect -666 532 5714 536
rect -666 528 -182 532
rect -682 394 6130 464
rect -680 -380 -476 394
rect 302 152 6130 394
rect 302 -380 532 152
rect 850 -380 1006 152
rect 1334 -380 1420 152
rect 1754 146 6130 152
rect 1754 144 3578 146
rect 1754 -380 1960 144
rect 2284 -380 2586 144
rect 2914 -380 2986 144
rect 3314 -380 3542 144
rect 3868 132 5136 146
rect 3868 -380 4162 132
rect 4494 -380 4590 132
rect 4906 -380 5136 132
rect 5460 -380 6130 146
rect -680 -594 6130 -380
rect -680 -775 6124 -594
rect -680 -881 -324 -775
rect -146 -881 6124 -775
rect -680 -954 6124 -881
<< viali >>
rect -493 1418 -387 1452
rect -324 -881 -146 -775
<< metal1 >>
rect -1006 1452 -106 1488
rect -1006 1418 -493 1452
rect -387 1418 -106 1452
rect 3354 1442 3402 1444
rect 3338 1440 4102 1442
rect 4692 1440 5860 1448
rect 2252 1438 5860 1440
rect 534 1436 562 1438
rect 1614 1436 5860 1438
rect -1006 1372 -106 1418
rect 92 1406 5860 1436
rect 92 1288 128 1406
rect 92 1282 126 1288
rect -38 1214 30 1222
rect -296 1196 -236 1206
rect -38 1196 -29 1214
rect -296 1194 -29 1196
rect -326 1164 -29 1194
rect -326 1148 -236 1164
rect -38 1162 -29 1164
rect 23 1162 30 1214
rect -38 1154 30 1162
rect -326 1086 -292 1148
rect 94 1118 126 1282
rect 178 1198 424 1244
rect -244 1082 128 1118
rect -328 642 -292 932
rect 178 756 212 1198
rect 534 1162 562 1406
rect 1614 1404 2314 1406
rect 3338 1404 5860 1406
rect 954 1264 1018 1270
rect 954 1212 960 1264
rect 1012 1260 1018 1264
rect 1012 1214 1108 1260
rect 1358 1214 1534 1268
rect 1012 1212 1018 1214
rect 954 1206 1018 1212
rect 462 1126 562 1162
rect 372 892 408 966
rect 1052 918 1088 996
rect 1140 956 1186 996
rect 1140 922 1174 956
rect 1202 922 1266 928
rect 1140 920 1266 922
rect 1038 912 1102 918
rect 356 886 420 892
rect 356 834 362 886
rect 414 834 420 886
rect 1038 860 1044 912
rect 1096 860 1102 912
rect 1140 888 1208 920
rect 1142 870 1208 888
rect 1202 868 1208 870
rect 1260 868 1266 920
rect 1202 860 1266 868
rect 1038 854 1102 860
rect 356 828 420 834
rect 178 720 678 756
rect -430 560 -400 562
rect -328 560 -290 642
rect -430 518 -288 560
rect -430 138 -400 518
rect -352 374 -286 380
rect -352 322 -344 374
rect -292 322 -286 374
rect -352 316 -286 322
rect -352 262 -322 316
rect -352 232 -274 262
rect 80 214 172 266
rect 80 174 120 214
rect -434 104 -298 138
rect -240 124 120 174
rect 80 112 120 124
rect 516 121 580 128
rect 516 69 522 121
rect 574 96 580 121
rect 574 69 582 96
rect 516 62 582 69
rect 554 -6 582 62
rect 644 34 674 720
rect 1046 109 1126 122
rect 1046 57 1061 109
rect 1113 80 1126 109
rect 1113 76 1184 80
rect 1358 76 1410 1214
rect 1616 1194 1646 1404
rect 2086 1264 2150 1270
rect 2086 1212 2092 1264
rect 2144 1256 2150 1264
rect 2144 1254 2198 1256
rect 2144 1212 2218 1254
rect 2086 1206 2218 1212
rect 1616 1174 1648 1194
rect 2274 1174 2314 1404
rect 3158 1268 3226 1274
rect 2760 1208 2874 1256
rect 3158 1216 3166 1268
rect 3218 1260 3226 1268
rect 3218 1224 3312 1260
rect 3218 1216 3226 1224
rect 3158 1210 3226 1216
rect 3354 1182 3402 1404
rect 3828 1236 3954 1268
rect 1564 1138 1648 1174
rect 2232 1130 2316 1174
rect 3316 1132 3406 1182
rect 1460 914 1500 988
rect 1446 906 1514 914
rect 1446 854 1453 906
rect 1505 854 1514 906
rect 1446 848 1514 854
rect 2142 146 2174 1040
rect 2820 894 2854 984
rect 2906 956 3264 994
rect 2552 860 2856 894
rect 2552 858 2854 860
rect 2552 168 2604 858
rect 2820 856 2854 858
rect 2544 162 2608 168
rect 1992 116 2176 146
rect 1113 57 1410 76
rect 1046 46 1410 57
rect 1108 42 1410 46
rect 1174 26 1410 42
rect 1452 76 1552 86
rect 1452 40 1602 76
rect 554 -34 668 -6
rect 74 -420 118 -160
rect 162 -284 206 -162
rect 716 -260 758 -176
rect 1104 -246 1148 -166
rect 1086 -254 1160 -246
rect 690 -275 776 -260
rect 690 -284 707 -275
rect 162 -327 707 -284
rect 759 -327 776 -275
rect 1086 -306 1097 -254
rect 1149 -306 1160 -254
rect 1086 -316 1160 -306
rect 162 -328 776 -327
rect 690 -342 776 -328
rect 1200 -344 1234 -192
rect 1270 -335 1336 -326
rect 1270 -344 1277 -335
rect 1200 -372 1277 -344
rect 1270 -387 1277 -372
rect 1329 -387 1336 -335
rect 1270 -394 1336 -387
rect 1452 -420 1480 40
rect 1518 18 1602 40
rect 1992 -14 2020 116
rect 2544 110 2550 162
rect 2602 110 2608 162
rect 2544 104 2608 110
rect 2552 102 2604 104
rect 2190 84 2264 90
rect 2190 72 2200 84
rect 2114 32 2200 72
rect 2252 32 2264 84
rect 3224 68 3288 74
rect 3224 62 3230 68
rect 2114 26 2264 32
rect 2614 24 2756 60
rect 3140 24 3230 62
rect 1510 -46 1574 -40
rect 1992 -44 2094 -14
rect 1510 -98 1516 -46
rect 1568 -98 1574 -46
rect 1510 -104 1574 -98
rect 1606 -258 1652 -196
rect 2142 -250 2188 -182
rect 1600 -264 1664 -258
rect 1600 -316 1606 -264
rect 1658 -316 1664 -264
rect 1600 -324 1664 -316
rect 2126 -264 2208 -250
rect 2126 -316 2141 -264
rect 2193 -316 2208 -264
rect 2126 -330 2208 -316
rect 2508 -420 2572 -418
rect 2614 -420 2642 24
rect 3224 16 3230 24
rect 3282 16 3288 68
rect 3828 56 3858 1236
rect 4050 1182 4092 1404
rect 4692 1402 5860 1404
rect 4000 1144 4092 1182
rect 4502 1234 4650 1270
rect 3900 930 3934 996
rect 3900 924 3968 930
rect 3900 906 3910 924
rect 3904 872 3910 906
rect 3962 872 3968 924
rect 3904 864 3968 872
rect 4502 626 4534 1234
rect 4716 1186 4748 1402
rect 4910 1302 4974 1308
rect 4910 1250 4916 1302
rect 4968 1294 4974 1302
rect 4968 1250 5044 1294
rect 5562 1268 5746 1270
rect 4910 1246 5044 1250
rect 4910 1242 4974 1246
rect 5540 1232 5746 1268
rect 4666 1146 4750 1186
rect 4574 932 4612 994
rect 4568 925 4634 932
rect 4568 873 4575 925
rect 4627 873 4634 925
rect 4568 866 4634 873
rect 4502 262 4536 626
rect 4990 412 5024 1002
rect 5092 998 5118 1006
rect 5076 936 5118 998
rect 5076 930 5140 936
rect 5076 878 5082 930
rect 5134 878 5140 930
rect 5076 872 5140 878
rect 5540 414 5582 1232
rect 5816 1184 5858 1402
rect 5764 1172 5858 1184
rect 5758 1108 5858 1172
rect 5758 1102 5848 1108
rect 5476 412 5582 414
rect 4990 392 5582 412
rect 5664 402 5700 1024
rect 4990 340 5494 392
rect 5546 340 5582 392
rect 4990 336 5582 340
rect 4204 67 4276 80
rect 3224 10 3288 16
rect 3412 52 3446 56
rect 3722 52 3860 56
rect 3412 14 3860 52
rect 4204 15 4214 67
rect 4266 58 4276 67
rect 4266 48 4342 58
rect 4500 48 4538 262
rect 4266 28 4538 48
rect 4616 48 4708 50
rect 4266 15 4536 28
rect 2686 -260 2724 -206
rect 2778 -238 3134 -198
rect 3184 -248 3226 -182
rect 3174 -254 3244 -248
rect 2672 -266 2738 -260
rect 2672 -318 2679 -266
rect 2731 -294 2738 -266
rect 2731 -318 2742 -294
rect 3174 -306 3183 -254
rect 3235 -306 3244 -254
rect 3174 -312 3244 -306
rect 2672 -324 2742 -318
rect 74 -422 1242 -420
rect 1366 -422 2642 -420
rect 74 -460 2642 -422
rect 74 -466 1490 -460
rect 1454 -468 1490 -466
rect -798 -744 -262 -742
rect -798 -775 338 -744
rect -798 -881 -324 -775
rect -146 -881 338 -775
rect 2508 -750 2572 -460
rect 2690 -476 2742 -324
rect 3412 -476 3446 14
rect 4204 6 4536 15
rect 4616 16 4756 48
rect 4204 2 4342 6
rect 4236 0 4342 2
rect 3580 -30 3662 -20
rect 3564 -36 3662 -30
rect 3564 -88 3570 -36
rect 3622 -42 3662 -36
rect 3622 -88 3666 -42
rect 3564 -94 3666 -88
rect 4228 -182 4292 -174
rect 3730 -256 3764 -208
rect 4228 -234 4234 -182
rect 4286 -234 4292 -182
rect 4228 -240 4292 -234
rect 3724 -263 3796 -256
rect 3724 -315 3732 -263
rect 3784 -315 3796 -263
rect 3724 -324 3796 -315
rect 4354 -270 4388 -224
rect 4354 -274 4424 -270
rect 4354 -280 4432 -274
rect 4354 -316 4370 -280
rect 4360 -332 4370 -316
rect 4422 -332 4432 -280
rect 4360 -338 4432 -332
rect 2688 -528 3446 -476
rect 3412 -532 3446 -528
rect 4616 -750 4650 16
rect 4776 -177 4842 -170
rect 4686 -278 4720 -228
rect 4776 -229 4782 -177
rect 4834 -229 4842 -177
rect 4776 -236 4842 -229
rect 4990 -278 5024 336
rect 5476 322 5582 336
rect 5476 312 5564 322
rect 5668 200 5700 402
rect 5164 148 5704 200
rect 5164 -24 5206 148
rect 5364 77 5428 86
rect 5364 68 5368 77
rect 5318 25 5368 68
rect 5420 25 5428 77
rect 5318 24 5428 25
rect 5364 18 5428 24
rect 5164 -56 5274 -24
rect 5166 -64 5274 -56
rect 4686 -306 5024 -278
rect 5324 -242 5366 -174
rect 5324 -253 5414 -242
rect 5324 -286 5351 -253
rect 5340 -305 5351 -286
rect 5403 -305 5414 -253
rect 5340 -314 5414 -305
rect 2508 -816 4650 -750
rect 2508 -818 4644 -816
rect 4506 -820 4644 -818
rect -798 -912 338 -881
rect -798 -914 -262 -912
<< rmetal1 >>
rect 2720 1256 2786 1276
rect 2720 1208 2760 1256
<< via1 >>
rect -29 1162 23 1214
rect 960 1212 1012 1264
rect 362 834 414 886
rect 1044 860 1096 912
rect 1208 868 1260 920
rect -344 322 -292 374
rect 522 69 574 121
rect 1061 57 1113 109
rect 2092 1212 2144 1264
rect 3166 1216 3218 1268
rect 1453 854 1505 906
rect 707 -327 759 -275
rect 1097 -306 1149 -254
rect 1277 -387 1329 -335
rect 2550 110 2602 162
rect 2200 32 2252 84
rect 1516 -98 1568 -46
rect 1606 -316 1658 -264
rect 2141 -316 2193 -264
rect 3230 16 3282 68
rect 3910 872 3962 924
rect 4916 1250 4968 1302
rect 4575 873 4627 925
rect 5082 878 5134 930
rect 5494 340 5546 392
rect 4214 15 4266 67
rect 2679 -318 2731 -266
rect 3183 -306 3235 -254
rect 3570 -88 3622 -36
rect 4234 -234 4286 -182
rect 3732 -315 3784 -263
rect 4370 -332 4422 -280
rect 4782 -229 4834 -177
rect 5368 25 5420 77
rect 5351 -305 5403 -253
<< metal2 >>
rect 970 1380 1002 1382
rect -18 1378 1002 1380
rect -18 1348 4948 1378
rect -18 1338 1002 1348
rect -18 1222 28 1338
rect 970 1270 1002 1338
rect 2732 1276 2762 1348
rect 4920 1308 4948 1348
rect 4910 1302 4974 1308
rect 954 1264 1018 1270
rect -38 1214 30 1222
rect -38 1162 -29 1214
rect 23 1162 30 1214
rect 954 1212 960 1264
rect 1012 1212 1018 1264
rect 2086 1264 2150 1270
rect 2086 1256 2092 1264
rect 1956 1212 2092 1256
rect 2144 1212 2150 1264
rect 954 1206 1018 1212
rect -38 1154 30 1162
rect 1202 920 1498 926
rect 1038 912 1102 918
rect 356 886 420 892
rect 356 834 362 886
rect 414 868 420 886
rect 414 838 734 868
rect 1038 860 1044 912
rect 1096 860 1102 912
rect 1202 868 1208 920
rect 1260 914 1498 920
rect 1260 906 1514 914
rect 1260 868 1453 906
rect 1202 866 1453 868
rect 1038 854 1102 860
rect 414 834 420 838
rect 356 828 420 834
rect 530 576 558 578
rect 706 576 734 838
rect 1052 582 1102 854
rect 1446 854 1453 866
rect 1505 854 1514 906
rect 1446 848 1514 854
rect 530 542 736 576
rect 530 540 592 542
rect -352 376 -286 380
rect -730 374 -286 376
rect -730 322 -344 374
rect -292 322 -286 374
rect -352 316 -286 322
rect 530 266 558 540
rect 1052 534 1706 582
rect 1052 530 1540 534
rect 530 234 1098 266
rect 530 128 558 234
rect 516 121 580 128
rect 1068 122 1098 234
rect 1666 256 1706 534
rect 1958 256 2012 1212
rect 2086 1206 2150 1212
rect 2720 1208 2786 1276
rect 3158 1268 3226 1274
rect 3158 1216 3166 1268
rect 3218 1216 3226 1268
rect 4910 1250 4916 1302
rect 4968 1250 4974 1302
rect 4910 1242 4974 1250
rect 3158 1210 3226 1216
rect 3162 256 3190 1210
rect 3904 924 3968 930
rect 3904 872 3910 924
rect 3962 872 3968 924
rect 3904 864 3968 872
rect 4568 925 4634 932
rect 4568 873 4575 925
rect 4627 916 4634 925
rect 5076 930 5140 936
rect 5076 916 5082 930
rect 4627 886 5082 916
rect 4627 873 4634 886
rect 4568 866 4634 873
rect 5076 878 5082 886
rect 5134 878 5140 930
rect 5076 872 5140 878
rect 1666 244 3190 256
rect 1666 212 3278 244
rect 3916 218 3956 864
rect 5544 414 5578 416
rect 5476 392 5578 414
rect 5476 340 5494 392
rect 5546 340 5578 392
rect 5476 338 5578 340
rect 5376 286 5582 338
rect 3912 216 4200 218
rect 3580 214 3674 216
rect 3912 214 4220 216
rect 516 69 522 121
rect 574 69 580 121
rect 516 62 580 69
rect 1046 109 1126 122
rect 1046 57 1061 109
rect 1113 57 1126 109
rect 1046 46 1126 57
rect 1510 -46 1574 -40
rect 1510 -98 1516 -46
rect 1568 -48 1574 -46
rect 1666 -48 1706 212
rect 2206 210 3170 212
rect 2206 90 2238 210
rect 2544 162 2608 168
rect 2544 110 2550 162
rect 2602 110 2608 162
rect 2544 104 2608 110
rect 2190 84 2264 90
rect 2190 32 2200 84
rect 2252 32 2264 84
rect 2190 26 2264 32
rect 1568 -82 1706 -48
rect 1568 -98 1574 -82
rect 1510 -104 1574 -98
rect 1086 -254 1664 -246
rect 690 -275 776 -260
rect 690 -327 707 -275
rect 759 -327 776 -275
rect 1086 -306 1097 -254
rect 1149 -264 1664 -254
rect 1149 -288 1606 -264
rect 1149 -306 1158 -288
rect 1086 -316 1158 -306
rect 1600 -316 1606 -288
rect 1658 -316 1664 -264
rect 1600 -324 1664 -316
rect 2126 -264 2208 -250
rect 2126 -316 2141 -264
rect 2193 -316 2208 -264
rect 2550 -278 2580 104
rect 3244 74 3276 212
rect 3580 180 4222 214
rect 3580 178 3674 180
rect 4164 178 4222 180
rect 3224 68 3288 74
rect 3224 16 3230 68
rect 3282 16 3288 68
rect 3224 10 3288 16
rect 3580 -30 3610 178
rect 4182 80 4222 178
rect 5376 86 5420 286
rect 4182 67 4276 80
rect 4182 15 4214 67
rect 4266 15 4276 67
rect 5364 77 5428 86
rect 5364 25 5368 77
rect 5420 25 5428 77
rect 5364 18 5428 25
rect 4182 2 4276 15
rect 4182 -4 4222 2
rect 3564 -36 3630 -30
rect 3564 -88 3570 -36
rect 3622 -88 3630 -36
rect 3564 -94 3630 -88
rect 4776 -174 4842 -170
rect 4228 -177 4842 -174
rect 4228 -182 4782 -177
rect 4228 -234 4234 -182
rect 4286 -224 4782 -182
rect 4286 -234 4292 -224
rect 4228 -240 4292 -234
rect 4776 -229 4782 -224
rect 4834 -229 4842 -177
rect 4776 -236 4842 -229
rect 3174 -254 3244 -248
rect 2672 -266 2738 -260
rect 2672 -278 2679 -266
rect 2550 -312 2679 -278
rect 690 -342 776 -327
rect 1270 -335 1336 -326
rect 2126 -330 2208 -316
rect 2672 -318 2679 -312
rect 2731 -318 2738 -266
rect 3174 -306 3183 -254
rect 3235 -306 3244 -254
rect 5340 -253 5414 -242
rect 3174 -312 3244 -306
rect 3724 -263 3796 -256
rect 2672 -324 2738 -318
rect 704 -634 760 -342
rect 1270 -387 1277 -335
rect 1329 -387 1336 -335
rect 1270 -394 1336 -387
rect 1284 -632 1334 -394
rect 2144 -632 2186 -330
rect 1282 -634 2188 -632
rect 700 -638 2188 -634
rect 3194 -638 3240 -312
rect 3724 -315 3732 -263
rect 3784 -315 3796 -263
rect 3724 -324 3796 -315
rect 4360 -280 4432 -274
rect 700 -644 3242 -638
rect 3732 -644 3786 -324
rect 4360 -332 4370 -280
rect 4422 -332 4432 -280
rect 5340 -305 5351 -253
rect 5403 -305 5414 -253
rect 5340 -314 5414 -305
rect 4360 -338 4432 -332
rect 700 -648 3786 -644
rect 4368 -648 4418 -338
rect 700 -650 4418 -648
rect 5348 -650 5396 -314
rect 700 -692 5396 -650
rect 1282 -700 5396 -692
rect 2056 -702 5396 -700
rect 3164 -704 5370 -702
rect 3164 -706 4410 -704
rect 3164 -708 3786 -706
rect 3732 -710 3786 -708
use sky130_fd_pr__nfet_01v8_KW5RPL  XM1
timestamp 1745430816
transform 1 0 -265 0 1 -14
box -201 -400 201 400
use sky130_fd_pr__nfet_01v8_KW5RPL  XM2
timestamp 1745430816
transform 1 0 141 0 1 -16
box -201 -400 201 400
use sky130_fd_pr__pfet_01v8_KBS6X7  XM3
timestamp 1745430816
transform 1 0 -267 0 1 1013
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM4
timestamp 1745430816
transform 1 0 689 0 1 -106
box -201 -300 201 300
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1745430816
transform 1 0 435 0 1 1059
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM11
timestamp 1745430816
transform 1 0 1173 0 1 -108
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_SFU2NW  XM12
timestamp 1745430816
transform 1 0 1585 0 1 -110
box -201 -300 201 300
use sky130_fd_pr__pfet_01v8_KBS6X7  XM13
timestamp 1745430816
transform 1 0 1113 0 1 1073
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM14
timestamp 1745430816
transform 1 0 1523 0 1 1073
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM19
timestamp 1745430816
transform 1 0 2203 0 1 1069
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM20
timestamp 1745430816
transform 1 0 2117 0 1 -116
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_SFU2NW  XM21
timestamp 1745430816
transform 1 0 3155 0 1 -120
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_SFU2NW  XM22
timestamp 1745430816
transform 1 0 2749 0 1 -120
box -201 -300 201 300
use sky130_fd_pr__pfet_01v8_KBS6X7  XM23
timestamp 1745430816
transform 1 0 2881 0 1 1067
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM24
timestamp 1745430816
transform 1 0 3285 0 1 1071
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM25
timestamp 1745430816
transform 1 0 3961 0 1 1081
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM26
timestamp 1745430816
transform 1 0 3703 0 1 -120
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_SFU2NW  XM27
timestamp 1745430816
transform 1 0 4327 0 1 -134
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_SFU2NW  XM28
timestamp 1745430816
transform 1 0 4747 0 1 -134
box -201 -300 201 300
use sky130_fd_pr__pfet_01v8_KBS6X7  XM29
timestamp 1745430816
transform 1 0 5049 0 1 1089
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM30
timestamp 1745430816
transform 1 0 4637 0 1 1083
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM31
timestamp 1745430816
transform 1 0 5731 0 1 1083
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM32
timestamp 1745430816
transform 1 0 5301 0 1 -114
box -201 -300 201 300
<< end >>
