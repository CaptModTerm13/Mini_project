magic
tech sky130A
magscale 1 2
timestamp 1745253145
<< locali >>
rect -6 524 28 536
rect 1324 -804 1392 -792
rect 842 -824 916 -812
rect 842 -858 868 -824
rect 902 -858 916 -824
rect 842 -868 916 -858
rect 1324 -860 1332 -804
rect 1382 -860 1392 -804
rect 1324 -868 1392 -860
rect 3448 -962 3548 -942
rect 3448 -1008 3460 -962
rect 3542 -1008 3548 -962
rect 3448 -1016 3548 -1008
rect 158 -1026 218 -1020
rect 158 -1064 164 -1026
rect 202 -1064 218 -1026
rect 158 -1068 218 -1064
<< viali >>
rect 2116 478 2152 516
rect 6306 486 6340 520
rect 4212 294 4270 362
rect 5718 -122 5762 -82
rect 3688 -222 3748 -174
rect 610 -334 656 -300
rect 1346 -326 1394 -290
rect 612 -336 652 -334
rect 2120 -436 2154 -390
rect 2942 -454 2994 -420
rect 3980 -472 4026 -424
rect 5226 -446 5264 -404
rect 6364 -466 6418 -414
rect 7404 -516 7442 -482
rect -542 -696 -490 -660
rect 868 -858 902 -824
rect 1332 -860 1382 -804
rect 2418 -1004 2546 -912
rect 3460 -1008 3542 -962
rect 4668 -972 4708 -936
rect 5712 -1008 5768 -950
rect -158 -1066 -120 -1028
rect 164 -1064 202 -1026
rect 6846 -1034 6886 -994
<< metal1 >>
rect 514 748 622 754
rect 2920 748 3012 756
rect -278 732 366 734
rect 514 732 526 748
rect -278 678 526 732
rect 610 732 622 748
rect 2100 740 2160 748
rect 2920 740 4112 748
rect 2100 732 4112 740
rect 610 690 4112 732
rect 610 682 3028 690
rect 610 678 2176 682
rect -278 658 366 678
rect 514 666 622 678
rect 1926 644 2020 650
rect 1926 622 1932 644
rect 26 614 1932 622
rect -6 574 30 612
rect 78 574 1932 614
rect -6 566 86 574
rect 1926 572 1932 574
rect 2010 572 2020 644
rect 1926 566 2020 572
rect -6 524 30 566
rect 82 534 518 536
rect 82 526 1732 534
rect 82 518 1752 526
rect 82 492 1690 518
rect 82 486 518 492
rect 1686 464 1690 492
rect 1746 464 1752 518
rect 1686 454 1752 464
rect 1936 404 1994 566
rect 2100 556 2160 678
rect 2100 522 2172 556
rect 2090 516 2172 522
rect 2090 478 2116 516
rect 2152 500 2172 516
rect 2152 478 2168 500
rect 2090 460 2168 478
rect 1936 394 2030 404
rect 2920 400 3012 682
rect 3972 654 4038 690
rect 5214 658 5280 682
rect 6294 658 7446 660
rect 5208 654 7446 658
rect 3972 608 7446 654
rect 3972 606 4992 608
rect -6 132 28 378
rect 1936 360 1994 394
rect 2020 354 2030 394
rect 1970 348 2030 354
rect 2026 276 2074 308
rect -586 78 28 132
rect 538 198 642 208
rect 538 124 540 198
rect 628 182 642 198
rect 1386 188 1794 222
rect 1386 186 1450 188
rect 628 124 654 182
rect 538 112 654 124
rect -584 -118 -550 78
rect -346 -34 -98 -32
rect -404 -46 -98 -34
rect -378 -86 -98 -46
rect -346 -88 -98 -86
rect -584 -162 -424 -118
rect 598 -228 654 112
rect 1386 48 1420 186
rect 1632 150 1710 160
rect 1494 148 1710 150
rect 1494 132 1642 148
rect 1480 120 1642 132
rect 1494 96 1642 120
rect 1694 96 1710 148
rect 1494 92 1710 96
rect 1494 82 1684 92
rect 1480 76 1538 82
rect 1634 80 1684 82
rect 1386 22 1480 48
rect 1386 14 1486 22
rect 1440 -16 1486 14
rect 1750 -110 1794 188
rect 2926 148 3006 400
rect 3972 358 4038 606
rect 5208 604 6348 608
rect 4354 390 4456 396
rect 4194 362 4284 376
rect 4194 358 4212 362
rect 3972 294 4212 358
rect 4270 294 4284 362
rect 4354 336 4362 390
rect 4450 336 4456 390
rect 4354 330 4456 336
rect 3514 282 3622 288
rect 3514 212 3520 282
rect 3612 212 3622 282
rect 3514 204 3622 212
rect 2026 138 2070 146
rect 2900 138 3054 148
rect 1936 -16 1978 134
rect 2020 82 2104 138
rect 2020 74 2108 82
rect 2020 72 2034 74
rect 2026 12 2034 72
rect 2096 38 2108 74
rect 2096 12 2104 38
rect 2026 2 2104 12
rect 2900 2 2908 138
rect 3040 2 3054 138
rect 2900 -8 3054 2
rect 3444 46 3544 52
rect 1936 -108 1980 -16
rect 1934 -110 2392 -108
rect 1442 -156 1488 -132
rect 1534 -156 1576 -140
rect 1750 -152 2392 -110
rect 1934 -154 2392 -152
rect 1534 -158 1578 -156
rect 1440 -202 1510 -196
rect 1540 -202 1578 -158
rect 598 -260 656 -228
rect 1440 -254 1446 -202
rect 1504 -230 1578 -202
rect 2208 -210 2272 -208
rect 2208 -214 2296 -210
rect 1504 -254 1510 -230
rect 1440 -260 1510 -254
rect 602 -294 656 -260
rect 2208 -266 2222 -214
rect 2286 -266 2296 -214
rect 2208 -274 2296 -266
rect 1332 -290 1404 -274
rect 2208 -276 2272 -274
rect 2176 -280 2272 -276
rect 1332 -294 1346 -290
rect 602 -300 666 -294
rect 602 -334 610 -300
rect 656 -334 666 -300
rect 602 -336 612 -334
rect 652 -336 666 -334
rect 602 -344 666 -336
rect 604 -352 666 -344
rect 1330 -326 1346 -294
rect 1394 -326 1404 -290
rect 2116 -304 2272 -280
rect 2116 -308 2206 -304
rect 1330 -340 1404 -326
rect -8 -400 54 -392
rect 738 -396 814 -390
rect -46 -402 54 -400
rect -46 -442 2 -402
rect 50 -442 54 -402
rect -46 -446 54 -442
rect 538 -398 990 -396
rect -46 -474 2 -446
rect 538 -450 748 -398
rect 802 -450 990 -398
rect 538 -462 990 -450
rect -380 -554 4 -474
rect 1330 -526 1392 -340
rect 2112 -390 2162 -308
rect 2112 -420 2120 -390
rect 2106 -436 2120 -420
rect 2154 -420 2162 -390
rect 2154 -436 2170 -420
rect 2106 -448 2170 -436
rect 1476 -498 1538 -492
rect 1476 -500 1598 -498
rect 1528 -504 1598 -500
rect 1984 -504 2044 -500
rect 1528 -506 2044 -504
rect -560 -660 -420 -652
rect -560 -696 -542 -660
rect -490 -696 -420 -660
rect -560 -718 -420 -696
rect -558 -1004 -422 -718
rect 456 -742 490 -692
rect 710 -726 814 -714
rect 710 -742 730 -726
rect 456 -784 730 -742
rect 710 -802 730 -784
rect 796 -742 814 -726
rect 946 -742 986 -676
rect 1330 -686 1380 -526
rect 1528 -542 1998 -506
rect 1476 -546 1998 -542
rect 1476 -548 1538 -546
rect 1408 -584 1488 -578
rect 1408 -646 1416 -584
rect 1482 -646 1488 -584
rect 1408 -652 1488 -646
rect 796 -784 986 -742
rect 796 -802 814 -784
rect 846 -822 928 -814
rect -558 -1028 -100 -1004
rect -558 -1066 -158 -1028
rect -120 -1066 -100 -1028
rect -558 -1076 -100 -1066
rect -558 -1266 -422 -1076
rect -44 -1118 -2 -842
rect 48 -932 96 -874
rect 846 -894 852 -822
rect 920 -894 928 -822
rect 846 -902 928 -894
rect 1036 -914 1078 -686
rect 1330 -792 1392 -686
rect 1324 -804 1392 -792
rect 1324 -860 1332 -804
rect 1382 -860 1392 -804
rect 1324 -868 1392 -860
rect 1328 -872 1392 -868
rect 1010 -922 1090 -914
rect 1010 -930 1020 -922
rect 578 -932 1020 -930
rect 48 -974 1020 -932
rect 578 -976 1020 -974
rect 1010 -984 1020 -976
rect 1084 -984 1090 -922
rect 1010 -992 1090 -984
rect 158 -1022 218 -1020
rect 550 -1022 636 -1008
rect 848 -1012 940 -1006
rect 848 -1022 856 -1012
rect 150 -1024 856 -1022
rect 150 -1026 560 -1024
rect 150 -1064 164 -1026
rect 202 -1064 560 -1026
rect 150 -1080 560 -1064
rect 630 -1080 856 -1024
rect 150 -1082 856 -1080
rect 926 -1024 940 -1012
rect 1328 -1024 1388 -872
rect 1524 -916 1578 -756
rect 1518 -922 1586 -916
rect 1518 -976 1524 -922
rect 1580 -976 1586 -922
rect 1518 -982 1586 -976
rect 926 -1082 1392 -1024
rect 1502 -1028 1598 -1022
rect 848 -1086 940 -1082
rect 1502 -1084 1508 -1028
rect 1592 -1084 1598 -1028
rect 1502 -1090 1598 -1084
rect -54 -1126 744 -1118
rect 1602 -1126 1692 -1124
rect -54 -1128 1692 -1126
rect -54 -1174 1616 -1128
rect -42 -1180 1616 -1174
rect 1674 -1180 1692 -1128
rect -42 -1184 1692 -1180
rect -42 -1190 1424 -1184
rect 1602 -1188 1692 -1184
rect 1734 -1272 1794 -546
rect 1966 -550 1998 -546
rect 2350 -524 2392 -154
rect 2926 -420 3006 -8
rect 3444 -20 3452 46
rect 3536 -20 3544 46
rect 3444 -26 3544 -20
rect 3590 -90 3640 -20
rect 3972 -54 4048 294
rect 4194 284 4284 294
rect 4286 116 4386 122
rect 4286 60 4296 116
rect 4378 60 4386 116
rect 4286 52 4386 60
rect 3488 -94 3640 -90
rect 3484 -116 3640 -94
rect 3484 -140 3636 -116
rect 3484 -402 3542 -140
rect 3678 -168 3764 -158
rect 3678 -228 3684 -168
rect 3756 -228 3764 -168
rect 3678 -236 3764 -228
rect 2926 -454 2942 -420
rect 2994 -454 3006 -420
rect 2926 -462 3006 -454
rect 2930 -466 3006 -462
rect 3466 -410 3566 -402
rect 3466 -470 3472 -410
rect 3556 -470 3566 -410
rect 3960 -424 4048 -54
rect 4242 -308 4330 -284
rect 4236 -314 4330 -308
rect 4236 -370 4242 -314
rect 4304 -362 4330 -314
rect 4304 -370 4312 -362
rect 4236 -376 4312 -370
rect 3960 -444 3980 -424
rect 3466 -476 3566 -470
rect 3968 -472 3980 -444
rect 4026 -444 4048 -424
rect 4428 -438 4462 118
rect 5214 -180 5280 604
rect 6298 528 6348 604
rect 6292 520 6356 528
rect 6292 486 6306 520
rect 6340 486 6356 520
rect 6292 476 6356 486
rect 6408 466 6502 474
rect 6408 396 6414 466
rect 6494 396 6502 466
rect 6408 388 6502 396
rect 5852 382 5946 388
rect 5852 322 5858 382
rect 5938 322 5946 382
rect 5852 314 5946 322
rect 5830 -28 5874 148
rect 5920 76 6008 86
rect 5920 10 5926 76
rect 5996 10 6008 76
rect 5920 4 6008 10
rect 6130 -6 6222 6
rect 6130 -28 6138 -6
rect 5830 -48 6138 -28
rect 5710 -82 5778 -68
rect 5832 -74 6138 -48
rect 5710 -90 5718 -82
rect 5762 -90 5778 -82
rect 5710 -142 5716 -90
rect 5770 -142 5778 -90
rect 6130 -88 6138 -74
rect 6208 -28 6222 -6
rect 6386 -28 6436 182
rect 6208 -74 6436 -28
rect 6208 -88 6222 -74
rect 6386 -82 6436 -74
rect 6130 -98 6222 -88
rect 6480 -92 6514 174
rect 6480 -114 6646 -92
rect 6482 -120 6646 -114
rect 6568 -124 6646 -120
rect 5710 -144 5778 -142
rect 5210 -196 5280 -180
rect 5210 -256 6424 -196
rect 5214 -388 5280 -256
rect 5426 -298 5508 -288
rect 5426 -358 5436 -298
rect 5498 -358 5508 -298
rect 5426 -366 5508 -358
rect 5214 -404 5282 -388
rect 4026 -472 4044 -444
rect 3968 -476 4044 -472
rect 3972 -482 4044 -476
rect 1966 -556 2046 -550
rect 1984 -560 2014 -556
rect 2350 -568 2636 -524
rect 2670 -568 3072 -518
rect 3352 -538 3604 -516
rect 3198 -572 3288 -542
rect 2128 -578 2176 -576
rect 1890 -636 1896 -584
rect 1952 -590 1958 -584
rect 2128 -590 2206 -578
rect 3198 -590 3218 -572
rect 1952 -636 1996 -590
rect 1890 -642 1996 -636
rect 2044 -640 2140 -590
rect 1896 -660 1996 -642
rect 2132 -644 2140 -640
rect 2202 -644 2206 -590
rect 2132 -650 2206 -644
rect 2696 -662 2722 -620
rect 3118 -624 3218 -590
rect 3276 -624 3288 -572
rect 3118 -634 3288 -624
rect 3198 -636 3288 -634
rect 3348 -572 3604 -538
rect 3640 -564 4100 -522
rect 2700 -740 2786 -732
rect 1952 -806 1998 -764
rect 2046 -804 2082 -786
rect 2590 -854 2630 -796
rect 2700 -808 2710 -740
rect 2778 -808 2786 -740
rect 2700 -818 2786 -808
rect 3028 -854 3068 -784
rect 2590 -856 3068 -854
rect 3348 -856 3416 -572
rect 4244 -596 4310 -590
rect 4244 -604 4252 -596
rect 3486 -612 3584 -606
rect 3486 -676 3492 -612
rect 3576 -676 3584 -612
rect 4158 -640 4252 -604
rect 4244 -648 4252 -640
rect 4304 -648 4310 -596
rect 4244 -652 4310 -648
rect 3486 -682 3584 -676
rect 2590 -892 3416 -856
rect 3028 -896 3068 -892
rect 2390 -912 2560 -900
rect 2390 -994 2418 -912
rect 2404 -1004 2418 -994
rect 2546 -1004 2560 -912
rect 2404 -1018 2560 -1004
rect 3438 -954 3564 -928
rect 3438 -1006 3452 -954
rect 3534 -962 3564 -954
rect 3438 -1008 3456 -1006
rect 3542 -1008 3564 -962
rect 3438 -1014 3564 -1008
rect 2694 -1042 2730 -1038
rect 2662 -1056 2758 -1042
rect 3650 -1052 3682 -778
rect 4064 -846 4100 -784
rect 4430 -808 4460 -438
rect 5214 -446 5226 -404
rect 5264 -446 5282 -404
rect 5214 -452 5282 -446
rect 4762 -508 4824 -504
rect 4762 -510 4850 -508
rect 4758 -564 4764 -510
rect 4818 -538 5378 -510
rect 4818 -564 4824 -538
rect 4758 -568 4824 -564
rect 4844 -568 5378 -538
rect 5460 -552 5496 -366
rect 6364 -404 6418 -256
rect 6454 -302 6558 -276
rect 6454 -360 6470 -302
rect 6536 -360 6558 -302
rect 6454 -376 6558 -360
rect 6352 -414 6436 -404
rect 6352 -466 6364 -414
rect 6418 -466 6436 -414
rect 6352 -474 6436 -466
rect 5614 -536 5848 -530
rect 5886 -536 6384 -526
rect 5614 -538 5858 -536
rect 4762 -570 4824 -568
rect 5460 -574 5502 -552
rect 5468 -616 5502 -574
rect 5406 -640 5502 -616
rect 5604 -580 5858 -538
rect 5406 -652 5500 -640
rect 4776 -778 4818 -774
rect 4740 -804 4818 -778
rect 4432 -846 4460 -808
rect 4064 -872 4460 -846
rect 4066 -880 4460 -872
rect 4432 -884 4460 -880
rect 4720 -810 4818 -804
rect 4720 -884 4728 -810
rect 4812 -884 4818 -810
rect 4720 -894 4818 -884
rect 4338 -918 4428 -912
rect 4338 -988 4346 -918
rect 4416 -928 4428 -918
rect 4664 -928 4720 -924
rect 4416 -936 4720 -928
rect 4416 -972 4668 -936
rect 4708 -972 4720 -936
rect 4416 -978 4720 -972
rect 4416 -988 4428 -978
rect 4664 -986 4720 -978
rect 4338 -996 4428 -988
rect 4868 -1052 4914 -790
rect 5304 -794 5322 -790
rect 5336 -794 5352 -784
rect 5304 -828 5352 -794
rect 5268 -834 5352 -828
rect 5268 -890 5278 -834
rect 5344 -838 5352 -834
rect 5604 -838 5656 -580
rect 5876 -584 6384 -536
rect 6480 -608 6518 -376
rect 5740 -620 5844 -614
rect 5740 -692 5748 -620
rect 5836 -692 5844 -620
rect 6430 -672 6518 -608
rect 6430 -674 6514 -672
rect 5740 -700 5844 -692
rect 5892 -824 5940 -782
rect 5344 -882 5656 -838
rect 5344 -890 5350 -882
rect 5604 -884 5656 -882
rect 5268 -896 5350 -890
rect 5698 -948 5782 -932
rect 5698 -1010 5712 -948
rect 5770 -1010 5782 -948
rect 5698 -1020 5782 -1010
rect 3646 -1054 4930 -1052
rect 5898 -1054 5940 -824
rect 6330 -866 6366 -794
rect 6612 -866 6646 -124
rect 7174 -104 7296 -84
rect 7174 -184 7192 -104
rect 7286 -132 7296 -104
rect 7286 -184 7300 -132
rect 7174 -204 7300 -184
rect 7222 -562 7300 -204
rect 7404 -474 7446 608
rect 7606 -284 7724 -272
rect 7606 -380 7614 -284
rect 7716 -380 7724 -284
rect 7606 -390 7724 -380
rect 7394 -482 7458 -474
rect 7394 -484 7404 -482
rect 7390 -516 7404 -484
rect 7442 -510 7458 -482
rect 7442 -516 7456 -510
rect 7390 -526 7456 -516
rect 6998 -620 7544 -562
rect 7658 -660 7696 -390
rect 7582 -710 7704 -660
rect 6872 -794 6946 -786
rect 6872 -846 6878 -794
rect 6930 -846 6946 -794
rect 6872 -852 6946 -846
rect 6330 -900 6648 -866
rect 6834 -984 6902 -980
rect 6834 -1042 6840 -984
rect 6894 -1042 6902 -984
rect 6834 -1048 6902 -1042
rect 3646 -1056 5940 -1054
rect 2662 -1060 5940 -1056
rect 2662 -1112 2678 -1060
rect 2736 -1096 5940 -1060
rect 2736 -1112 2766 -1096
rect 3646 -1098 5940 -1096
rect 4868 -1100 4914 -1098
rect 2662 -1126 2766 -1112
rect 2662 -1128 2758 -1126
rect 2232 -1138 2338 -1132
rect 2232 -1210 2238 -1138
rect 2330 -1152 2338 -1138
rect 3252 -1142 3412 -1126
rect 3252 -1152 3268 -1142
rect 2330 -1158 2632 -1152
rect 2788 -1158 3268 -1152
rect 2330 -1210 3268 -1158
rect 2232 -1218 3268 -1210
rect 2284 -1220 3268 -1218
rect 2632 -1230 2788 -1220
rect 1734 -1338 1738 -1272
rect 1790 -1338 1794 -1272
rect 3252 -1262 3268 -1220
rect 3396 -1262 3412 -1142
rect 5894 -1236 5940 -1098
rect 3252 -1282 3412 -1262
rect 5896 -1256 5940 -1236
rect 7018 -1256 7064 -840
rect 7448 -844 7524 -834
rect 7448 -900 7454 -844
rect 7516 -900 7524 -844
rect 7448 -908 7524 -900
rect 5896 -1292 7064 -1256
rect 5896 -1298 7058 -1292
rect 5896 -1300 5940 -1298
rect 1734 -1366 1794 -1338
<< via1 >>
rect 526 678 610 748
rect 1932 572 2010 644
rect 1690 464 1746 518
rect 540 124 628 198
rect 1642 96 1694 148
rect 4362 336 4450 390
rect 3520 212 3612 282
rect 2034 12 2096 74
rect 2908 2 3040 138
rect 1446 -254 1504 -202
rect 2222 -266 2286 -214
rect 748 -450 802 -398
rect 730 -802 796 -726
rect 1416 -646 1482 -584
rect 852 -824 920 -822
rect 852 -858 868 -824
rect 868 -858 902 -824
rect 902 -858 920 -824
rect 852 -894 920 -858
rect 1020 -984 1084 -922
rect 560 -1080 630 -1024
rect 856 -1082 926 -1012
rect 1524 -976 1580 -922
rect 1508 -1084 1592 -1028
rect 1616 -1180 1674 -1128
rect 3452 -20 3536 46
rect 4296 60 4378 116
rect 3684 -174 3756 -168
rect 3684 -222 3688 -174
rect 3688 -222 3748 -174
rect 3748 -222 3756 -174
rect 3684 -228 3756 -222
rect 3472 -470 3556 -410
rect 4242 -370 4304 -314
rect 6414 396 6494 466
rect 5858 322 5938 382
rect 5926 10 5996 76
rect 5716 -122 5718 -90
rect 5718 -122 5762 -90
rect 5762 -122 5770 -90
rect 5716 -142 5770 -122
rect 6138 -88 6208 -6
rect 5436 -358 5498 -298
rect 1896 -636 1952 -584
rect 2140 -644 2202 -590
rect 3218 -624 3276 -572
rect 2710 -808 2778 -740
rect 3492 -676 3576 -612
rect 4252 -648 4304 -596
rect 2418 -1004 2546 -912
rect 3452 -962 3534 -954
rect 3452 -1006 3460 -962
rect 3456 -1008 3460 -1006
rect 3460 -1008 3534 -962
rect 4764 -564 4818 -510
rect 6470 -360 6536 -302
rect 4728 -884 4812 -810
rect 4346 -988 4416 -918
rect 5278 -890 5344 -834
rect 5748 -692 5836 -620
rect 5712 -950 5770 -948
rect 5712 -1008 5768 -950
rect 5768 -1008 5770 -950
rect 5712 -1010 5770 -1008
rect 7192 -184 7286 -104
rect 7614 -380 7716 -284
rect 6878 -846 6930 -794
rect 6840 -994 6894 -984
rect 6840 -1034 6846 -994
rect 6846 -1034 6886 -994
rect 6886 -1034 6894 -994
rect 6840 -1042 6894 -1034
rect 2678 -1112 2736 -1060
rect 2238 -1210 2330 -1138
rect 1738 -1338 1790 -1272
rect 3268 -1262 3396 -1142
rect 7454 -900 7516 -844
<< metal2 >>
rect 7902 1206 8042 1286
rect 750 1148 8194 1206
rect 744 1104 8194 1148
rect 514 748 622 754
rect 514 678 526 748
rect 610 678 622 748
rect 744 712 802 1104
rect 6426 740 6478 742
rect 514 666 622 678
rect 548 208 620 666
rect 538 198 642 208
rect 538 124 540 198
rect 628 124 642 198
rect 538 112 642 124
rect 746 -390 794 712
rect 5554 696 6484 740
rect 5550 670 6484 696
rect 4380 654 4416 656
rect 3476 650 4416 654
rect 1926 644 4416 650
rect 1926 572 1932 644
rect 2010 606 4416 644
rect 2010 602 3500 606
rect 2010 572 2020 602
rect 1926 566 2020 572
rect 1674 518 1754 534
rect 1674 464 1690 518
rect 1746 464 1754 518
rect 1674 400 1754 464
rect 2072 400 2166 402
rect 1674 384 2166 400
rect 4380 396 4416 606
rect 5550 396 5618 670
rect 6426 474 6478 670
rect 6408 466 6502 474
rect 6408 396 6414 466
rect 6494 396 6502 466
rect 1678 352 2166 384
rect 4354 390 5646 396
rect 1632 148 1710 160
rect 1632 96 1642 148
rect 1694 96 1710 148
rect 2126 124 2164 352
rect 4354 336 4362 390
rect 4450 336 5646 390
rect 4354 330 5646 336
rect 5848 382 5950 392
rect 6408 388 6502 396
rect 5848 322 5858 382
rect 5938 322 5950 382
rect 5848 312 5950 322
rect 3504 288 3632 296
rect 3504 204 3514 288
rect 3622 204 3632 288
rect 3504 194 3632 204
rect 2900 138 3054 148
rect 2126 118 2178 124
rect 1632 92 1710 96
rect 1634 80 1694 92
rect 1636 78 1694 80
rect 1636 50 1690 78
rect 1616 -184 1690 50
rect 2026 74 2104 84
rect 2026 12 2034 74
rect 2096 12 2104 74
rect 2026 2 2104 12
rect 2038 -176 2090 2
rect 2136 -30 2178 118
rect 2900 106 2908 138
rect 2236 26 2908 106
rect 1906 -178 2098 -176
rect 1440 -202 1510 -196
rect 1440 -254 1446 -202
rect 1504 -254 1510 -202
rect 1440 -260 1510 -254
rect 738 -398 814 -390
rect 738 -450 748 -398
rect 802 -450 814 -398
rect 738 -456 814 -450
rect 1444 -578 1478 -260
rect 1408 -584 1488 -578
rect 1408 -646 1416 -584
rect 1482 -646 1488 -584
rect 1408 -652 1488 -646
rect 722 -802 730 -726
rect 796 -802 802 -726
rect 730 -986 796 -802
rect 846 -822 928 -814
rect 846 -894 852 -822
rect 920 -894 928 -822
rect 846 -902 928 -894
rect 550 -1024 636 -1008
rect 550 -1042 560 -1024
rect 558 -1080 560 -1042
rect 630 -1042 636 -1024
rect 558 -1276 630 -1080
rect 730 -1094 800 -986
rect 856 -1006 912 -902
rect 1010 -922 1090 -914
rect 1010 -984 1020 -922
rect 1084 -932 1090 -922
rect 1518 -922 1586 -916
rect 1518 -932 1524 -922
rect 1084 -976 1524 -932
rect 1580 -976 1586 -922
rect 1084 -984 1090 -976
rect 1010 -992 1090 -984
rect 1022 -996 1084 -992
rect 848 -1012 940 -1006
rect 848 -1082 856 -1012
rect 926 -1082 940 -1012
rect 1518 -1022 1586 -976
rect 1618 -998 1688 -184
rect 1898 -230 2098 -178
rect 1898 -584 1940 -230
rect 2126 -312 2164 -30
rect 2236 -204 2304 26
rect 2900 2 2908 26
rect 3040 2 3054 138
rect 4286 116 4386 122
rect 4286 60 4296 116
rect 4378 60 4386 116
rect 4286 52 4386 60
rect 5920 76 6008 86
rect 2900 -8 3054 2
rect 3444 46 3544 52
rect 3444 -20 3452 46
rect 3536 -20 3544 46
rect 3444 -26 3544 -20
rect 3454 -62 3496 -26
rect 4330 -60 4368 52
rect 5920 10 5926 76
rect 5996 10 6008 76
rect 5920 4 6008 10
rect 4330 -62 4370 -60
rect 3454 -76 4370 -62
rect 3456 -106 4370 -76
rect 4330 -118 4370 -106
rect 5710 -90 5778 -88
rect 4330 -122 4788 -118
rect 4330 -158 4790 -122
rect 5710 -136 5716 -90
rect 2226 -210 2304 -204
rect 2212 -214 2304 -210
rect 2212 -266 2222 -214
rect 2286 -250 2304 -214
rect 3678 -168 3764 -158
rect 3678 -228 3684 -168
rect 3756 -188 3764 -168
rect 4356 -188 4404 -186
rect 3756 -228 4404 -188
rect 3678 -236 3764 -228
rect 4356 -250 4404 -228
rect 2286 -266 2300 -250
rect 2212 -274 2296 -266
rect 4242 -294 4330 -284
rect 4242 -308 4252 -294
rect 4236 -312 4252 -308
rect 2126 -316 2826 -312
rect 3180 -314 4252 -312
rect 3180 -316 4242 -314
rect 2126 -362 4242 -316
rect 4320 -352 4330 -294
rect 2126 -578 2164 -362
rect 2748 -364 4242 -362
rect 3180 -370 4242 -364
rect 4304 -362 4330 -352
rect 4304 -370 4312 -362
rect 3182 -542 3226 -370
rect 4236 -376 4312 -370
rect 3466 -410 3566 -402
rect 3466 -470 3472 -410
rect 3556 -470 3566 -410
rect 3466 -476 3566 -470
rect 3182 -572 3288 -542
rect 1890 -636 1896 -584
rect 1952 -636 1958 -584
rect 2126 -590 2206 -578
rect 2126 -610 2140 -590
rect 1890 -642 1958 -636
rect 2132 -644 2140 -610
rect 2202 -644 2206 -590
rect 3182 -592 3218 -572
rect 3198 -624 3218 -592
rect 3276 -624 3288 -572
rect 3500 -606 3530 -476
rect 4246 -550 4308 -376
rect 4364 -410 4404 -250
rect 4244 -596 4310 -550
rect 3198 -636 3288 -624
rect 3486 -612 3584 -606
rect 2132 -650 2206 -644
rect 3486 -676 3492 -612
rect 3576 -676 3584 -612
rect 4244 -648 4252 -596
rect 4304 -648 4310 -596
rect 4244 -652 4310 -648
rect 3486 -682 3584 -676
rect 2700 -740 2786 -732
rect 2700 -808 2710 -740
rect 2778 -808 2786 -740
rect 2700 -818 2786 -808
rect 2404 -912 2560 -900
rect 2404 -940 2418 -912
rect 848 -1086 940 -1082
rect 1502 -1028 1594 -1022
rect 1502 -1084 1508 -1028
rect 1592 -1084 1594 -1028
rect 856 -1088 914 -1086
rect 1502 -1090 1518 -1084
rect 734 -1254 800 -1094
rect 1508 -1098 1518 -1090
rect 1580 -1090 1594 -1084
rect 1580 -1098 1590 -1090
rect 1508 -1106 1574 -1098
rect 1622 -1122 1688 -998
rect 1618 -1124 1688 -1122
rect 2386 -1004 2418 -940
rect 2546 -1004 2560 -912
rect 2386 -1018 2560 -1004
rect 1602 -1128 1692 -1124
rect 1602 -1180 1616 -1128
rect 1674 -1134 1692 -1128
rect 2232 -1134 2338 -1132
rect 1674 -1138 2338 -1134
rect 1674 -1180 2238 -1138
rect 1602 -1188 2238 -1180
rect 1610 -1198 2238 -1188
rect 2232 -1210 2238 -1198
rect 2330 -1210 2338 -1138
rect 2232 -1218 2338 -1210
rect 730 -1272 1822 -1254
rect 550 -1414 632 -1276
rect 730 -1338 1738 -1272
rect 1790 -1338 1822 -1272
rect 730 -1360 1822 -1338
rect 2386 -1410 2504 -1018
rect 2714 -1036 2762 -818
rect 4356 -912 4404 -410
rect 4752 -504 4790 -158
rect 5598 -142 5716 -136
rect 5770 -142 5778 -90
rect 5598 -170 5760 -142
rect 5426 -298 5508 -288
rect 5426 -358 5436 -298
rect 5498 -358 5508 -298
rect 5426 -366 5508 -358
rect 4752 -510 4824 -504
rect 4752 -558 4764 -510
rect 4758 -564 4764 -558
rect 4818 -564 4824 -510
rect 4758 -568 4824 -564
rect 4762 -570 4824 -568
rect 4720 -810 4818 -804
rect 4720 -884 4728 -810
rect 4812 -854 4818 -810
rect 5268 -834 5350 -828
rect 5268 -854 5278 -834
rect 4812 -884 5278 -854
rect 4720 -888 5278 -884
rect 4720 -894 4818 -888
rect 5268 -890 5278 -888
rect 5344 -890 5350 -834
rect 5268 -896 5350 -890
rect 4338 -918 4428 -912
rect 3446 -954 3544 -948
rect 3446 -1006 3452 -954
rect 3446 -1008 3456 -1006
rect 3534 -1008 3544 -954
rect 4338 -988 4346 -918
rect 4416 -988 4428 -918
rect 4338 -996 4428 -988
rect 3446 -1014 3544 -1008
rect 2662 -1052 2764 -1036
rect 2662 -1118 2672 -1052
rect 2744 -1118 2764 -1052
rect 2662 -1124 2764 -1118
rect 2662 -1128 2758 -1124
rect 3252 -1136 3412 -1126
rect 3252 -1268 3260 -1136
rect 3404 -1268 3412 -1136
rect 3252 -1282 3412 -1268
rect 3452 -1140 3532 -1014
rect 4356 -1032 4396 -996
rect 4360 -1140 4396 -1032
rect 3452 -1142 4396 -1140
rect 5598 -1142 5642 -170
rect 5752 -300 5822 -296
rect 5942 -300 5996 4
rect 6130 -6 6222 6
rect 6130 -88 6138 -6
rect 6208 -88 6222 -6
rect 6130 -98 6222 -88
rect 6148 -134 6200 -98
rect 7174 -104 7296 -84
rect 7174 -126 7192 -104
rect 6736 -134 7192 -126
rect 6146 -176 7192 -134
rect 6736 -178 7192 -176
rect 7174 -184 7192 -178
rect 7286 -184 7296 -104
rect 7174 -204 7296 -184
rect 6454 -294 6558 -276
rect 5752 -346 5998 -300
rect 5752 -614 5786 -346
rect 6454 -366 6464 -294
rect 6540 -366 6558 -294
rect 6454 -376 6558 -366
rect 7606 -284 7724 -272
rect 7606 -380 7614 -284
rect 7716 -286 7724 -284
rect 7718 -376 7724 -286
rect 7716 -380 7724 -376
rect 7606 -390 7724 -380
rect 5740 -620 5844 -614
rect 5740 -692 5748 -620
rect 5836 -692 5844 -620
rect 5740 -700 5844 -692
rect 6872 -794 6946 -786
rect 6872 -846 6878 -794
rect 6930 -846 6946 -794
rect 6872 -852 6946 -846
rect 7448 -844 7524 -834
rect 6880 -892 6928 -852
rect 7234 -892 7290 -888
rect 7448 -892 7454 -844
rect 6880 -900 7454 -892
rect 7516 -900 7524 -844
rect 6880 -908 7524 -900
rect 7902 -866 8042 1104
rect 6880 -918 7510 -908
rect 6886 -924 7510 -918
rect 5702 -948 5780 -940
rect 5702 -1010 5712 -948
rect 5770 -1010 5780 -948
rect 5702 -1018 5780 -1010
rect 6834 -984 6902 -980
rect 3452 -1144 5676 -1142
rect 5718 -1144 5756 -1018
rect 6834 -1042 6840 -984
rect 6894 -1042 6902 -984
rect 6834 -1050 6902 -1042
rect 3452 -1146 5756 -1144
rect 6840 -1146 6886 -1050
rect 3452 -1182 6890 -1146
rect 3452 -1410 3532 -1182
rect 4306 -1188 6890 -1182
rect 4360 -1190 4396 -1188
rect 5656 -1192 6890 -1188
rect 5656 -1194 5742 -1192
rect 7234 -1210 7290 -924
rect 7902 -1210 8040 -866
rect 7234 -1290 8042 -1210
rect 7902 -1304 8040 -1290
rect 2386 -1414 3544 -1410
rect 550 -1452 3544 -1414
rect 554 -1508 3544 -1452
rect 2390 -1510 3544 -1508
<< via2 >>
rect 5858 322 5938 382
rect 3514 282 3622 288
rect 3514 212 3520 282
rect 3520 212 3612 282
rect 3612 212 3622 282
rect 3514 204 3622 212
rect 4252 -314 4320 -294
rect 4252 -352 4304 -314
rect 4304 -352 4320 -314
rect 1518 -1084 1580 -1042
rect 1518 -1098 1580 -1084
rect 5436 -358 5498 -298
rect 2672 -1060 2744 -1052
rect 2672 -1112 2678 -1060
rect 2678 -1112 2736 -1060
rect 2736 -1112 2744 -1060
rect 2672 -1118 2744 -1112
rect 3260 -1142 3404 -1136
rect 3260 -1262 3268 -1142
rect 3268 -1262 3396 -1142
rect 3396 -1262 3404 -1142
rect 3260 -1268 3404 -1262
rect 6464 -302 6540 -294
rect 6464 -360 6470 -302
rect 6470 -360 6536 -302
rect 6536 -360 6540 -302
rect 6464 -366 6540 -360
rect 7614 -376 7716 -286
rect 7716 -376 7718 -286
<< metal3 >>
rect 5862 570 5936 572
rect 3530 516 5936 570
rect 3526 496 5936 516
rect 3526 296 3622 496
rect 5862 392 5936 496
rect 5848 382 5950 392
rect 5848 322 5858 382
rect 5938 322 5950 382
rect 5848 312 5950 322
rect 5862 300 5936 312
rect 3504 288 3632 296
rect 3504 284 3514 288
rect 3322 212 3514 284
rect 1510 -1034 1586 -1032
rect 1510 -1036 1590 -1034
rect 1510 -1042 1880 -1036
rect 1508 -1098 1518 -1042
rect 1580 -1056 1880 -1042
rect 2662 -1052 2758 -1042
rect 2662 -1054 2672 -1052
rect 2638 -1056 2672 -1054
rect 1580 -1098 2672 -1056
rect 1508 -1106 1590 -1098
rect 1808 -1116 2672 -1098
rect 2662 -1118 2672 -1116
rect 2744 -1118 2758 -1052
rect 2662 -1128 2758 -1118
rect 3322 -1126 3386 212
rect 3504 204 3514 212
rect 3622 204 3632 288
rect 3504 194 3632 204
rect 4242 -294 4330 -284
rect 6454 -286 6558 -276
rect 7606 -286 7724 -272
rect 4242 -352 4252 -294
rect 4320 -298 4330 -294
rect 5426 -294 5508 -288
rect 6454 -294 7614 -286
rect 5426 -298 6464 -294
rect 4320 -352 5436 -298
rect 4242 -358 5436 -352
rect 5498 -358 6464 -298
rect 4242 -362 4330 -358
rect 5426 -366 5508 -358
rect 6454 -366 6464 -358
rect 6540 -366 7614 -294
rect 6454 -372 7614 -366
rect 6454 -376 6558 -372
rect 7606 -376 7614 -372
rect 7718 -376 7724 -286
rect 7606 -390 7724 -376
rect 3252 -1136 3412 -1126
rect 3252 -1268 3260 -1136
rect 3404 -1268 3412 -1136
rect 3252 -1282 3412 -1268
use sky130_fd_pr__nfet_01v8_KW5RPL  XM1
timestamp 1745227888
transform 1 0 -401 0 1 -318
box -211 -410 211 410
use sky130_fd_pr__nfet_01v8_KW5RPL  XM2
timestamp 1745227888
transform 1 0 23 0 1 -676
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_KBS6X7  XM3
timestamp 1745253145
transform 1 0 55 0 1 429
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM4
timestamp 1745227888
transform 1 0 1011 0 1 -594
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM5
timestamp 1745253145
transform 1 0 517 0 1 -595
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM11
timestamp 1745227888
transform 1 0 1505 0 1 -676
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM12
timestamp 1745227888
transform 1 0 1509 0 1 -54
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM13
timestamp 1745253145
transform 1 0 1999 0 1 211
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM14
timestamp 1745253145
transform 1 0 2017 0 1 -693
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM19
timestamp 1745253145
transform 1 0 3091 0 1 -701
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM20
timestamp 1745227888
transform 1 0 2653 0 1 -702
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM21
timestamp 1745227888
transform 1 0 3623 0 1 -706
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM22
timestamp 1745227888
transform 1 0 3561 0 1 76
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM23
timestamp 1745253145
transform 1 0 4399 0 1 189
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM24
timestamp 1745253145
transform 1 0 4123 0 1 -705
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM25
timestamp 1745253145
transform 1 0 5371 0 1 -703
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM26
timestamp 1745227888
transform 1 0 4841 0 1 -700
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM27
timestamp 1745227888
transform 1 0 5869 0 1 -714
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_SFU2NW  XM28
timestamp 1745227888
transform 1 0 5899 0 1 160
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_KBS6X7  XM29
timestamp 1745253145
transform 1 0 6451 0 1 245
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM30
timestamp 1745253145
transform 1 0 6391 0 1 -713
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_KBS6X7  XM31
timestamp 1745253145
transform 1 0 7547 0 1 -761
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_SFU2NW  XM32
timestamp 1745227888
transform 1 0 6993 0 1 -750
box -211 -310 211 310
<< end >>
