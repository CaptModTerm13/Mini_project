* Extracted by KLayout

* cell ros_ckt
* pin SUBSTRATE
.SUBCKT ros_ckt 21
* net 21 SUBSTRATE
* device instance $1 r0 *1 19.805,5.405 PMOS
M$1 20 3 11 24 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $2 r0 *1 14.405,5.335 PMOS
M$2 18 19 3 25 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $3 r0 *1 25.245,5.445 PMOS
M$3 17 13 5 23 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $4 r0 *1 28.655,5.415 PMOS
M$4 20 5 8 22 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $5 r0 *1 5.565,5.365 PMOS
M$5 16 13 6 27 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $6 r0 *1 16.425,5.355 PMOS
M$6 20 6 18 25 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $7 r0 *1 11.015,5.345 PMOS
M$7 20 6 10 26 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $8 r0 *1 23.185,5.415 PMOS
M$8 20 11 17 23 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $9 r0 *1 2.175,5.295 PMOS
M$9 20 15 12 28 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $10 r0 *1 7.615,5.365 PMOS
M$10 20 12 16 27 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $11 r0 *1 -1.335,5.065 PMOS
M$11 20 13 13 29 PMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $12 r0 *1 13.745,-0.6 NMOS
M$12 9 1 3 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $13 r0 *1 7.925,-0.55 NMOS
M$13 4 1 6 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $14 r0 *1 23.735,-0.67 NMOS
M$14 7 1 5 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $15 r0 *1 3.445,-0.53 NMOS
M$15 2 15 12 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $16 r0 *1 5.865,-0.54 NMOS
M$16 2 12 4 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $17 r0 *1 10.585,-0.58 NMOS
M$17 2 6 10 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $18 r0 *1 15.775,-0.6 NMOS
M$18 2 6 9 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $19 r0 *1 18.515,-0.6 NMOS
M$19 2 3 11 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $20 r0 *1 21.635,-0.67 NMOS
M$20 2 11 7 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $21 r0 *1 26.505,-0.57 NMOS
M$21 2 5 8 21 NMOS L=0.15U W=1U AS=0.29P AD=0.29P PS=2.58U PD=2.58U
* device instance $22 r0 *1 0.705,-0.08 NMOS
M$22 2 1 1 21 NMOS L=0.15U W=2U AS=0.58P AD=0.58P PS=4.58U PD=4.58U
* device instance $23 r0 *1 -1.325,-0.07 NMOS
M$23 1 14 13 21 NMOS L=0.15U W=2U AS=0.58P AD=0.58P PS=4.58U PD=4.58U
.ENDS ros_ckt
